module mem_exponent (clk, addr, cen, wen, data, q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;// Note
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b11000010111111000000000000000000 ;
        2:  q   <=  32'b11000010111110100000000000000000 ;
        3:  q   <=  32'b11000010111110000000000000000000 ;
        4:  q   <=  32'b11000010111101100000000000000000 ;
        5:  q   <=  32'b11000010111101000000000000000000 ;
        6:  q   <=  32'b11000010111100100000000000000000 ;
        7:  q   <=  32'b11000010111100000000000000000000 ;
        8:  q   <=  32'b11000010111011100000000000000000 ;
        9:  q   <=  32'b11000010111011000000000000000000 ;
        10:  q   <=  32'b11000010111010100000000000000000 ;
        11:  q   <=  32'b11000010111010000000000000000000 ;
        12:  q   <=  32'b11000010111001100000000000000000 ;
        13:  q   <=  32'b11000010111001000000000000000000 ;
        14:  q   <=  32'b11000010111000100000000000000000 ;
        15:  q   <=  32'b11000010111000000000000000000000 ;
        16:  q   <=  32'b11000010110111100000000000000000 ;
        17:  q   <=  32'b11000010110111000000000000000000 ;
        18:  q   <=  32'b11000010110110100000000000000000 ;
        19:  q   <=  32'b11000010110110000000000000000000 ;
        20:  q   <=  32'b11000010110101100000000000000000 ;
        21:  q   <=  32'b11000010110101000000000000000000 ;
        22:  q   <=  32'b11000010110100100000000000000000 ;
        23:  q   <=  32'b11000010110100000000000000000000 ;
        24:  q   <=  32'b11000010110011100000000000000000 ;
        25:  q   <=  32'b11000010110011000000000000000000 ;
        26:  q   <=  32'b11000010110010100000000000000000 ;
        27:  q   <=  32'b11000010110010000000000000000000 ;
        28:  q   <=  32'b11000010110001100000000000000000 ;
        29:  q   <=  32'b11000010110001000000000000000000 ;
        30:  q   <=  32'b11000010110000100000000000000000 ;
        31:  q   <=  32'b11000010110000000000000000000000 ;
        32:  q   <=  32'b11000010101111100000000000000000 ;
        33:  q   <=  32'b11000010101111000000000000000000 ;
        34:  q   <=  32'b11000010101110100000000000000000 ;
        35:  q   <=  32'b11000010101110000000000000000000 ;
        36:  q   <=  32'b11000010101101100000000000000000 ;
        37:  q   <=  32'b11000010101101000000000000000000 ;
        38:  q   <=  32'b11000010101100100000000000000000 ;
        39:  q   <=  32'b11000010101100000000000000000000 ;
        40:  q   <=  32'b11000010101011100000000000000000 ;
        41:  q   <=  32'b11000010101011000000000000000000 ;
        42:  q   <=  32'b11000010101010100000000000000000 ;
        43:  q   <=  32'b11000010101010000000000000000000 ;
        44:  q   <=  32'b11000010101001100000000000000000 ;
        45:  q   <=  32'b11000010101001000000000000000000 ;
        46:  q   <=  32'b11000010101000100000000000000000 ;
        47:  q   <=  32'b11000010101000000000000000000000 ;
        48:  q   <=  32'b11000010100111100000000000000000 ;
        49:  q   <=  32'b11000010100111000000000000000000 ;
        50:  q   <=  32'b11000010100110100000000000000000 ;
        51:  q   <=  32'b11000010100110000000000000000000 ;
        52:  q   <=  32'b11000010100101100000000000000000 ;
        53:  q   <=  32'b11000010100101000000000000000000 ;
        54:  q   <=  32'b11000010100100100000000000000000 ;
        55:  q   <=  32'b11000010100100000000000000000000 ;
        56:  q   <=  32'b11000010100011100000000000000000 ;
        57:  q   <=  32'b11000010100011000000000000000000 ;
        58:  q   <=  32'b11000010100010100000000000000000 ;
        59:  q   <=  32'b11000010100010000000000000000000 ;
        60:  q   <=  32'b11000010100001100000000000000000 ;
        61:  q   <=  32'b11000010100001000000000000000000 ;
        62:  q   <=  32'b11000010100000100000000000000000 ;
        63:  q   <=  32'b11000010100000000000000000000000 ;
        64:  q   <=  32'b11000010011111000000000000000000 ;
        65:  q   <=  32'b11000010011110000000000000000000 ;
        66:  q   <=  32'b11000010011101000000000000000000 ;
        67:  q   <=  32'b11000010011100000000000000000000 ;
        68:  q   <=  32'b11000010011011000000000000000000 ;
        69:  q   <=  32'b11000010011010000000000000000000 ;
        70:  q   <=  32'b11000010011001000000000000000000 ;
        71:  q   <=  32'b11000010011000000000000000000000 ;
        72:  q   <=  32'b11000010010111000000000000000000 ;
        73:  q   <=  32'b11000010010110000000000000000000 ;
        74:  q   <=  32'b11000010010101000000000000000000 ;
        75:  q   <=  32'b11000010010100000000000000000000 ;
        76:  q   <=  32'b11000010010011000000000000000000 ;
        77:  q   <=  32'b11000010010010000000000000000000 ;
        78:  q   <=  32'b11000010010001000000000000000000 ;
        79:  q   <=  32'b11000010010000000000000000000000 ;
        80:  q   <=  32'b11000010001111000000000000000000 ;
        81:  q   <=  32'b11000010001110000000000000000000 ;
        82:  q   <=  32'b11000010001101000000000000000000 ;
        83:  q   <=  32'b11000010001100000000000000000000 ;
        84:  q   <=  32'b11000010001011000000000000000000 ;
        85:  q   <=  32'b11000010001010000000000000000000 ;
        86:  q   <=  32'b11000010001001000000000000000000 ;
        87:  q   <=  32'b11000010001000000000000000000000 ;
        88:  q   <=  32'b11000010000111000000000000000000 ;
        89:  q   <=  32'b11000010000110000000000000000000 ;
        90:  q   <=  32'b11000010000101000000000000000000 ;
        91:  q   <=  32'b11000010000100000000000000000000 ;
        92:  q   <=  32'b11000010000011000000000000000000 ;
        93:  q   <=  32'b11000010000010000000000000000000 ;
        94:  q   <=  32'b11000010000001000000000000000000 ;
        95:  q   <=  32'b11000010000000000000000000000000 ;
        96:  q   <=  32'b11000001111110000000000000000000 ;
        97:  q   <=  32'b11000001111100000000000000000000 ;
        98:  q   <=  32'b11000001111010000000000000000000 ;
        99:  q   <=  32'b11000001111000000000000000000000 ;
        100:  q   <=  32'b11000001110110000000000000000000 ;
        101:  q   <=  32'b11000001110100000000000000000000 ;
        102:  q   <=  32'b11000001110010000000000000000000 ;
        103:  q   <=  32'b11000001110000000000000000000000 ;
        104:  q   <=  32'b11000001101110000000000000000000 ;
        105:  q   <=  32'b11000001101100000000000000000000 ;
        106:  q   <=  32'b11000001101010000000000000000000 ;
        107:  q   <=  32'b11000001101000000000000000000000 ;
        108:  q   <=  32'b11000001100110000000000000000000 ;
        109:  q   <=  32'b11000001100100000000000000000000 ;
        110:  q   <=  32'b11000001100010000000000000000000 ;
        111:  q   <=  32'b11000001100000000000000000000000 ;
        112:  q   <=  32'b11000001011100000000000000000000 ;
        113:  q   <=  32'b11000001011000000000000000000000 ;
        114:  q   <=  32'b11000001010100000000000000000000 ;
        115:  q   <=  32'b11000001010000000000000000000000 ;
        116:  q   <=  32'b11000001001100000000000000000000 ;
        117:  q   <=  32'b11000001001000000000000000000000 ;
        118:  q   <=  32'b11000001000100000000000000000000 ;
        119:  q   <=  32'b11000001000000000000000000000000 ;
        120:  q   <=  32'b11000000111000000000000000000000 ;
        121:  q   <=  32'b11000000110000000000000000000000 ;
        122:  q   <=  32'b11000000101000000000000000000000 ;
        123:  q   <=  32'b11000000100000000000000000000000 ;
        124:  q   <=  32'b11000000010000000000000000000000 ;
        125:  q   <=  32'b11000000000000000000000000000000 ;
        126:  q   <=  32'b10111111100000000000000000000000 ;
        127:  q   <=  32'b00000000000000000000000000000000 ;
        128:  q   <=  32'b00111111100000000000000000000000 ;
        129:  q   <=  32'b01000000000000000000000000000000 ;
        130:  q   <=  32'b01000000010000000000000000000000 ;
        131:  q   <=  32'b01000000100000000000000000000000 ;
        132:  q   <=  32'b01000000101000000000000000000000 ;
        133:  q   <=  32'b01000000110000000000000000000000 ;
        134:  q   <=  32'b01000000111000000000000000000000 ;
        135:  q   <=  32'b01000001000000000000000000000000 ;
        136:  q   <=  32'b01000001000100000000000000000000 ;
        137:  q   <=  32'b01000001001000000000000000000000 ;
        138:  q   <=  32'b01000001001100000000000000000000 ;
        139:  q   <=  32'b01000001010000000000000000000000 ;
        140:  q   <=  32'b01000001010100000000000000000000 ;
        141:  q   <=  32'b01000001011000000000000000000000 ;
        142:  q   <=  32'b01000001011100000000000000000000 ;
        143:  q   <=  32'b01000001100000000000000000000000 ;
        144:  q   <=  32'b01000001100010000000000000000000 ;
        145:  q   <=  32'b01000001100100000000000000000000 ;
        146:  q   <=  32'b01000001100110000000000000000000 ;
        147:  q   <=  32'b01000001101000000000000000000000 ;
        148:  q   <=  32'b01000001101010000000000000000000 ;
        149:  q   <=  32'b01000001101100000000000000000000 ;
        150:  q   <=  32'b01000001101110000000000000000000 ;
        151:  q   <=  32'b01000001110000000000000000000000 ;
        152:  q   <=  32'b01000001110010000000000000000000 ;
        153:  q   <=  32'b01000001110100000000000000000000 ;
        154:  q   <=  32'b01000001110110000000000000000000 ;
        155:  q   <=  32'b01000001111000000000000000000000 ;
        156:  q   <=  32'b01000001111010000000000000000000 ;
        157:  q   <=  32'b01000001111100000000000000000000 ;
        158:  q   <=  32'b01000001111110000000000000000000 ;
        159:  q   <=  32'b01000010000000000000000000000000 ;
        160:  q   <=  32'b01000010000001000000000000000000 ;
        161:  q   <=  32'b01000010000010000000000000000000 ;
        162:  q   <=  32'b01000010000011000000000000000000 ;
        163:  q   <=  32'b01000010000100000000000000000000 ;
        164:  q   <=  32'b01000010000101000000000000000000 ;
        165:  q   <=  32'b01000010000110000000000000000000 ;
        166:  q   <=  32'b01000010000111000000000000000000 ;
        167:  q   <=  32'b01000010001000000000000000000000 ;
        168:  q   <=  32'b01000010001001000000000000000000 ;
        169:  q   <=  32'b01000010001010000000000000000000 ;
        170:  q   <=  32'b01000010001011000000000000000000 ;
        171:  q   <=  32'b01000010001100000000000000000000 ;
        172:  q   <=  32'b01000010001101000000000000000000 ;
        173:  q   <=  32'b01000010001110000000000000000000 ;
        174:  q   <=  32'b01000010001111000000000000000000 ;
        175:  q   <=  32'b01000010010000000000000000000000 ;
        176:  q   <=  32'b01000010010001000000000000000000 ;
        177:  q   <=  32'b01000010010010000000000000000000 ;
        178:  q   <=  32'b01000010010011000000000000000000 ;
        179:  q   <=  32'b01000010010100000000000000000000 ;
        180:  q   <=  32'b01000010010101000000000000000000 ;
        181:  q   <=  32'b01000010010110000000000000000000 ;
        182:  q   <=  32'b01000010010111000000000000000000 ;
        183:  q   <=  32'b01000010011000000000000000000000 ;
        184:  q   <=  32'b01000010011001000000000000000000 ;
        185:  q   <=  32'b01000010011010000000000000000000 ;
        186:  q   <=  32'b01000010011011000000000000000000 ;
        187:  q   <=  32'b01000010011100000000000000000000 ;
        188:  q   <=  32'b01000010011101000000000000000000 ;
        189:  q   <=  32'b01000010011110000000000000000000 ;
        190:  q   <=  32'b01000010011111000000000000000000 ;
        191:  q   <=  32'b01000010100000000000000000000000 ;
        192:  q   <=  32'b01000010100000100000000000000000 ;
        193:  q   <=  32'b01000010100001000000000000000000 ;
        194:  q   <=  32'b01000010100001100000000000000000 ;
        195:  q   <=  32'b01000010100010000000000000000000 ;
        196:  q   <=  32'b01000010100010100000000000000000 ;
        197:  q   <=  32'b01000010100011000000000000000000 ;
        198:  q   <=  32'b01000010100011100000000000000000 ;
        199:  q   <=  32'b01000010100100000000000000000000 ;
        200:  q   <=  32'b01000010100100100000000000000000 ;
        201:  q   <=  32'b01000010100101000000000000000000 ;
        202:  q   <=  32'b01000010100101100000000000000000 ;
        203:  q   <=  32'b01000010100110000000000000000000 ;
        204:  q   <=  32'b01000010100110100000000000000000 ;
        205:  q   <=  32'b01000010100111000000000000000000 ;
        206:  q   <=  32'b01000010100111100000000000000000 ;
        207:  q   <=  32'b01000010101000000000000000000000 ;
        208:  q   <=  32'b01000010101000100000000000000000 ;
        209:  q   <=  32'b01000010101001000000000000000000 ;
        210:  q   <=  32'b01000010101001100000000000000000 ;
        211:  q   <=  32'b01000010101010000000000000000000 ;
        212:  q   <=  32'b01000010101010100000000000000000 ;
        213:  q   <=  32'b01000010101011000000000000000000 ;
        214:  q   <=  32'b01000010101011100000000000000000 ;
        215:  q   <=  32'b01000010101100000000000000000000 ;
        216:  q   <=  32'b01000010101100100000000000000000 ;
        217:  q   <=  32'b01000010101101000000000000000000 ;
        218:  q   <=  32'b01000010101101100000000000000000 ;
        219:  q   <=  32'b01000010101110000000000000000000 ;
        220:  q   <=  32'b01000010101110100000000000000000 ;
        221:  q   <=  32'b01000010101111000000000000000000 ;
        222:  q   <=  32'b01000010101111100000000000000000 ;
        223:  q   <=  32'b01000010110000000000000000000000 ;
        224:  q   <=  32'b01000010110000100000000000000000 ;
        225:  q   <=  32'b01000010110001000000000000000000 ;
        226:  q   <=  32'b01000010110001100000000000000000 ;
        227:  q   <=  32'b01000010110010000000000000000000 ;
        228:  q   <=  32'b01000010110010100000000000000000 ;
        229:  q   <=  32'b01000010110011000000000000000000 ;
        230:  q   <=  32'b01000010110011100000000000000000 ;
        231:  q   <=  32'b01000010110100000000000000000000 ;
        232:  q   <=  32'b01000010110100100000000000000000 ;
        233:  q   <=  32'b01000010110101000000000000000000 ;
        234:  q   <=  32'b01000010110101100000000000000000 ;
        235:  q   <=  32'b01000010110110000000000000000000 ;
        236:  q   <=  32'b01000010110110100000000000000000 ;
        237:  q   <=  32'b01000010110111000000000000000000 ;
        238:  q   <=  32'b01000010110111100000000000000000 ;
        239:  q   <=  32'b01000010111000000000000000000000 ;
        240:  q   <=  32'b01000010111000100000000000000000 ;
        241:  q   <=  32'b01000010111001000000000000000000 ;
        242:  q   <=  32'b01000010111001100000000000000000 ;
        243:  q   <=  32'b01000010111010000000000000000000 ;
        244:  q   <=  32'b01000010111010100000000000000000 ;
        245:  q   <=  32'b01000010111011000000000000000000 ;
        246:  q   <=  32'b01000010111011100000000000000000 ;
        247:  q   <=  32'b01000010111100000000000000000000 ;
        248:  q   <=  32'b01000010111100100000000000000000 ;
        249:  q   <=  32'b01000010111101000000000000000000 ;
        250:  q   <=  32'b01000010111101100000000000000000 ;
        251:  q   <=  32'b01000010111110000000000000000000 ;
        252:  q   <=  32'b01000010111110100000000000000000 ;
        253:  q   <=  32'b01000010111111000000000000000000 ;
        254:  q   <=  32'b01000010111111100000000000000000;
        default: q <= 0;
    endcase
end
endmodule
