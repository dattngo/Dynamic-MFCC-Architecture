module set_cofig (clk, 
