module mem_input_data (clk, addr, cen, wen, data, q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;// Note
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00111111000010011010010010001101 ;
        2:  q   <=  32'b00111111111010101011110010111110 ;
        3:  q   <=  32'b11000000000100001001000011110010 ;
        4:  q   <=  32'b00111111010111001011011101100100 ;
        5:  q   <=  32'b00111110101000110011010100110010 ;
        6:  q   <=  32'b10111111101001110110001001010100 ;
        7:  q   <=  32'b10111110110111011111111111000110 ;
        8:  q   <=  32'b00111110101011110110110001111001 ;
        9:  q   <=  32'b01000000011001010000010001110100 ;
        10:  q   <=  32'b01000000001100010011111001110100 ;
        11:  q   <=  32'b10111111101011001100100100011000 ;
        12:  q   <=  32'b01000000010000100011110000101111 ;
        13:  q   <=  32'b00111111001110011011010000010111 ;
        14:  q   <=  32'b10111101100000010010001011101001 ;
        15:  q   <=  32'b00111111001101101111100101100100 ;
        16:  q   <=  32'b10111110010100011110001010011111 ;
        17:  q   <=  32'b10111101111111100011111101100100 ;
        18:  q   <=  32'b00111111101111101010111001101001 ;
        19:  q   <=  32'b00111111101101000101101100111101 ;
        20:  q   <=  32'b00111111101101010110011010001111 ;
        21:  q   <=  32'b00111111001010111110011100111100 ;
        22:  q   <=  32'b10111111100110101000111011101110 ;
        23:  q   <=  32'b00111111001101111001110011110011 ;
        24:  q   <=  32'b00111111110100001010101110001100 ;
        25:  q   <=  32'b00111110111110100101000001001000 ;
        26:  q   <=  32'b00111111100001000111000011010010 ;
        27:  q   <=  32'b00111111001110100001010100100100 ;
        28:  q   <=  32'b10111110100110110101110010011011 ;
        29:  q   <=  32'b00111110100101100111011001010010 ;
        30:  q   <=  32'b10111111010010011000101101011101 ;
        31:  q   <=  32'b00111111011000110110110111100101 ;
        32:  q   <=  32'b10111111100100101101001100110001 ;
        33:  q   <=  32'b10111111100010001101000010111111 ;
        34:  q   <=  32'b10111111010011110011101101001110 ;
        35:  q   <=  32'b11000000001111000110111100100110 ;
        36:  q   <=  32'b00111111101110000001110011011000 ;
        37:  q   <=  32'b00111110101001100111111101011111 ;
        38:  q   <=  32'b10111111010000010100001011111011 ;
        39:  q   <=  32'b00111111101011110110010111110001 ;
        40:  q   <=  32'b10111111110110110001001011111000 ;
        41:  q   <=  32'b10111101110100010110010001111100 ;
        42:  q   <=  32'b10111110011101110011110111100100 ;
        43:  q   <=  32'b00111110101000110110111100010000 ;
        44:  q   <=  32'b00111110101000000010111100000000 ;
        45:  q   <=  32'b10111111010111010110100011000101 ;
        46:  q   <=  32'b10111100111101100010111000100010 ;
        47:  q   <=  32'b10111110001010001101011000001011 ;
        48:  q   <=  32'b00111111001000001011000101101100 ;
        49:  q   <=  32'b00111111100010111111000000100001 ;
        50:  q   <=  32'b00111111100011011111110010101010 ;
        51:  q   <=  32'b10111111010111010001100001011001 ;
        52:  q   <=  32'b00111101100111100110111001110001 ;
        53:  q   <=  32'b10111111100110110110100000101111 ;
        54:  q   <=  32'b10111111100011101000011100110001 ;
        55:  q   <=  32'b10111011111000000111000001010100 ;
        56:  q   <=  32'b00111111110001000010110100111010 ;
        57:  q   <=  32'b10111111010001010000100011010011 ;
        58:  q   <=  32'b00111110101111100010010101011101 ;
        59:  q   <=  32'b10111110011001101111111110011000 ;
        60:  q   <=  32'b00111111100011110000010110000110 ;
        61:  q   <=  32'b10111111100010110110011001110101 ;
        62:  q   <=  32'b00111101000001010101101011111001 ;
        63:  q   <=  32'b00111111000011010111001001101001 ;
        64:  q   <=  32'b00111111100011001110000011001011 ;
        65:  q   <=  32'b00111111110001011010100010111100 ;
        66:  q   <=  32'b00111101101011111111110010101001 ;
        67:  q   <=  32'b10111111101111101110110001101110 ;
        68:  q   <=  32'b10111111001111100000011101111110 ;
        69:  q   <=  32'b10111111100001111110000111101001 ;
        70:  q   <=  32'b01000000000101100110110111100100 ;
        71:  q   <=  32'b10111111000111011001100000010101 ;
        72:  q   <=  32'b00111111001111111000000111110101 ;
        73:  q   <=  32'b10111110010001010000100101011011 ;
        74:  q   <=  32'b00111111011000110111101111111001 ;
        75:  q   <=  32'b10111111010000111100110100101000 ;
        76:  q   <=  32'b10111111101100110111110110001100 ;
        77:  q   <=  32'b10111111101101100001000001101010 ;
        78:  q   <=  32'b00111110111110011111010010001101 ;
        79:  q   <=  32'b10111110001101011010000111010101 ;
        80:  q   <=  32'b10111110010010001100001000111110 ;
        81:  q   <=  32'b00111111101101011010101111110100 ;
        82:  q   <=  32'b00111110100101010100101010001100 ;
        83:  q   <=  32'b00111110010010101000111011111011 ;
        84:  q   <=  32'b00111111110010110011100110111001 ;
        85:  q   <=  32'b10111111010011011111000101111011 ;
        86:  q   <=  32'b00111111001100100101010111111010 ;
        87:  q   <=  32'b00111111010101011100100001010110 ;
        88:  q   <=  32'b10111110011110011001000001110110 ;
        89:  q   <=  32'b00111110010111001101100010011110 ;
        90:  q   <=  32'b10111111100101010011101001011111 ;
        91:  q   <=  32'b10111111100100101111000000011101 ;
        92:  q   <=  32'b00111101110101101100100010001110 ;
        93:  q   <=  32'b00111111001110001110010110100011 ;
        94:  q   <=  32'b01000000001001010111100010110000 ;
        95:  q   <=  32'b10111111001010101011100101011000 ;
        96:  q   <=  32'b00111110001111111101001110110100 ;
        97:  q   <=  32'b10111101101010001111001011010110 ;
        98:  q   <=  32'b10111111111101110110110101001011 ;
        99:  q   <=  32'b10111110111000001100000000101011 ;
        100:  q   <=  32'b10111111111001011011100000001001 ;
        101:  q   <=  32'b00111111010101110010001011011001 ;
        102:  q   <=  32'b10111111011000110101011000010010 ;
        103:  q   <=  32'b00111101110011001111110101111000 ;
        104:  q   <=  32'b10111111000010110110011000111111 ;
        105:  q   <=  32'b00111110100110110110011100010011 ;
        106:  q   <=  32'b10111111000110011010111100000000 ;
        107:  q   <=  32'b00111110111110101101110010111100 ;
        108:  q   <=  32'b00111111001111010100011011100110 ;
        109:  q   <=  32'b00111111110110110001111100100011 ;
        110:  q   <=  32'b10111110010001101100100001010001 ;
        111:  q   <=  32'b11000000000010001101101011010000 ;
        112:  q   <=  32'b10111111010101101110111101001001 ;
        113:  q   <=  32'b00111111101011010110001101011000 ;
        114:  q   <=  32'b10111111100010010011110001100010 ;
        115:  q   <=  32'b00111111011101100000000100010010 ;
        116:  q   <=  32'b00111101111111100000110111010010 ;
        117:  q   <=  32'b00111111101101111110010110101100 ;
        118:  q   <=  32'b10111111111110101111111011000101 ;
        119:  q   <=  32'b10111110010010100111000101100111 ;
        120:  q   <=  32'b10111111100110101001101010101110 ;
        121:  q   <=  32'b01000000001110100001110011001101 ;
        122:  q   <=  32'b00111111010100110100000110001011 ;
        123:  q   <=  32'b00111111101100001000001000100111 ;
        124:  q   <=  32'b10111111100001110111001001110011 ;
        125:  q   <=  32'b10111110111011111110111001100001 ;
        126:  q   <=  32'b10111110100010111000000100011100 ;
        127:  q   <=  32'b00111111100011001001100100101101 ;
        128:  q   <=  32'b10111110100011100100010100111010 ;
        129:  q   <=  32'b00111111001100111001100000111000 ;
        130:  q   <=  32'b11000000000000110101000011110101 ;
        131:  q   <=  32'b10111110101101010010101111010011 ;
        132:  q   <=  32'b10111111010100101101011010010001 ;
        133:  q   <=  32'b10111111110010011101110100000001 ;
        134:  q   <=  32'b00111111000000100000101010100000 ;
        135:  q   <=  32'b00111110100100000110000000110111 ;
        136:  q   <=  32'b00111101000010010010001000110011 ;
        137:  q   <=  32'b10111111101010101011010111110101 ;
        138:  q   <=  32'b00111111100100000101000110101010 ;
        139:  q   <=  32'b00111110101100110100101010110111 ;
        140:  q   <=  32'b10111110100110010001111100101110 ;
        141:  q   <=  32'b00111100101110111000001101011111 ;
        142:  q   <=  32'b10111110100001100010010001000100 ;
        143:  q   <=  32'b10111111111000000000011011110101 ;
        144:  q   <=  32'b10111110100100100100000011011000 ;
        145:  q   <=  32'b10111111010101001101010001101111 ;
        146:  q   <=  32'b10111111011110101010110101000011 ;
        147:  q   <=  32'b10111111100101000000010011111000 ;
        148:  q   <=  32'b10111111000010001001011100110010 ;
        149:  q   <=  32'b11000000000000000010101100101111 ;
        150:  q   <=  32'b00111111011101101101011110111101 ;
        151:  q   <=  32'b00111111000001010010001010101000 ;
        152:  q   <=  32'b10111100101001000001000101110010 ;
        153:  q   <=  32'b10111101000011100110110000100000 ;
        154:  q   <=  32'b10111111010011000101010001110010 ;
        155:  q   <=  32'b00111111100000100110010001000111 ;
        156:  q   <=  32'b10111110000010000110101000101001 ;
        157:  q   <=  32'b10111111001101101110101101110010 ;
        158:  q   <=  32'b00111111101011001111101000110101 ;
        159:  q   <=  32'b10111110011001100010101001100010 ;
        160:  q   <=  32'b10111111000101101100101010011011 ;
        161:  q   <=  32'b10111110100101100110011011011111 ;
        162:  q   <=  32'b10111111010110010001000110110001 ;
        163:  q   <=  32'b10111111100011110110000001011101 ;
        164:  q   <=  32'b01000000001000011010100111111010 ;
        165:  q   <=  32'b00111111110100111110011101011000 ;
        166:  q   <=  32'b00111110100111010111010100111111 ;
        167:  q   <=  32'b10111111101000001110100101000001 ;
        168:  q   <=  32'b10111111010111011000111101010000 ;
        169:  q   <=  32'b10111110001101001100010101011011 ;
        170:  q   <=  32'b00111111010010101001101000111110 ;
        171:  q   <=  32'b10111111101010100111111100011110 ;
        172:  q   <=  32'b11000000000101010001110010001011 ;
        173:  q   <=  32'b10111111101110010111110000000101 ;
        174:  q   <=  32'b00111110101010101100000111101110 ;
        175:  q   <=  32'b00111110110010000101111101111111 ;
        176:  q   <=  32'b00111110111001110100001010000110 ;
        177:  q   <=  32'b10111110000001010110100101010111 ;
        178:  q   <=  32'b00111110001111000001100011111110 ;
        179:  q   <=  32'b10111110111100111100101001010100 ;
        180:  q   <=  32'b00111111010111001010110101110010 ;
        181:  q   <=  32'b10111111101011100100110000000001 ;
        182:  q   <=  32'b00111110111010001111100110100010 ;
        183:  q   <=  32'b10111111010110010100010100000100 ;
        184:  q   <=  32'b10111110101010110111011001001101 ;
        185:  q   <=  32'b00111111000011011000001100110101 ;
        186:  q   <=  32'b00111111100001010000000011101100 ;
        187:  q   <=  32'b10111111100011110000111011001000 ;
        188:  q   <=  32'b00111111101000010101110101000011 ;
        189:  q   <=  32'b00111111001010001111111100100100 ;
        190:  q   <=  32'b10111101100010101111110100011000 ;
        191:  q   <=  32'b10111110010001111110100000010000 ;
        192:  q   <=  32'b10111110010111101101010000110010 ;
        193:  q   <=  32'b10111110100110110011000011101100 ;
        194:  q   <=  32'b00111100101111001100101000101101 ;
        195:  q   <=  32'b00111101010100100001010111010110 ;
        196:  q   <=  32'b00111111010100110111100011011001 ;
        197:  q   <=  32'b00111111110000110111001111111000 ;
        198:  q   <=  32'b00111110111011110000111101101000 ;
        199:  q   <=  32'b10111110010101101011111100010111 ;
        200:  q   <=  32'b00111111001000000000110001111001 ;
        201:  q   <=  32'b00111110001110111001111111101101 ;
        202:  q   <=  32'b10111111100000111100111101101100 ;
        203:  q   <=  32'b00111111011100110000000000110011 ;
        204:  q   <=  32'b00111110100111010011011100111000 ;
        205:  q   <=  32'b00111110000010100110101101001100 ;
        206:  q   <=  32'b00111111000000111110011100101111 ;
        207:  q   <=  32'b00111110100001011101011100001100 ;
        208:  q   <=  32'b10111111011100010000010100110110 ;
        209:  q   <=  32'b10111110001001100011101111011000 ;
        210:  q   <=  32'b10111110000101011000111101011000 ;
        211:  q   <=  32'b10111111000010000011000111100101 ;
        212:  q   <=  32'b00111111110101110100111100101011 ;
        213:  q   <=  32'b10111111011000000010111111001100 ;
        214:  q   <=  32'b10111110111101111011011010011011 ;
        215:  q   <=  32'b10111111001101100100010111101110 ;
        216:  q   <=  32'b10111111100101100100110010010110 ;
        217:  q   <=  32'b10111110010001001101101001101111 ;
        218:  q   <=  32'b10111110100011000101001011101110 ;
        219:  q   <=  32'b00111111110000111101100101101010 ;
        220:  q   <=  32'b10111110011111110000000001010111 ;
        221:  q   <=  32'b10111111100010000011100000100101 ;
        222:  q   <=  32'b00111111110011010011111000010110 ;
        223:  q   <=  32'b00111111100111100000100111110111 ;
        224:  q   <=  32'b10111110011010110010001100110010 ;
        225:  q   <=  32'b10111111110000001100100111010111 ;
        226:  q   <=  32'b10111110111000111010011001000001 ;
        227:  q   <=  32'b10111110000111111010111100000001 ;
        228:  q   <=  32'b00111110100011010101100011010001 ;
        229:  q   <=  32'b10111110100001011011011100111101 ;
        230:  q   <=  32'b00111110111000110000100000110010 ;
        231:  q   <=  32'b00111110110010001010011001011011 ;
        232:  q   <=  32'b10111111101000000001011000111111 ;
        233:  q   <=  32'b10111111011100101010110110010001 ;
        234:  q   <=  32'b10111111001111011011100100100001 ;
        235:  q   <=  32'b10111111000000100000000001010100 ;
        236:  q   <=  32'b10111110101001000010001001111001 ;
        237:  q   <=  32'b00111100010011000100101011110011 ;
        238:  q   <=  32'b11000000010000011101111000001010 ;
        239:  q   <=  32'b10111110111010011111110111010010 ;
        240:  q   <=  32'b00111111100111110000100010001100 ;
        241:  q   <=  32'b10111111100010001000100110101011 ;
        242:  q   <=  32'b00111111011011110000100011001111 ;
        243:  q   <=  32'b00111110101100110101110101000110 ;
        244:  q   <=  32'b10111100111011011001110101111110 ;
        245:  q   <=  32'b00111110001110101101010010111101 ;
        246:  q   <=  32'b10111111110010000101001111000001 ;
        247:  q   <=  32'b10111101101011010010001100001000 ;
        248:  q   <=  32'b00111111110011010100111000011101 ;
        249:  q   <=  32'b00111101110010010110101010001110 ;
        250:  q   <=  32'b00111101001010010111011101100000 ;
        251:  q   <=  32'b10111111001110111111001010000001 ;
        252:  q   <=  32'b10111100111111000110110100010011 ;
        253:  q   <=  32'b00111110011011011110110001100000 ;
        254:  q   <=  32'b00111110110110100100111101111000 ;
        255:  q   <=  32'b10111110101111101110000011001001 ;
        256:  q   <=  32'b10111110011100100010000100100110 ;
        257:  q   <=  32'b01000000000000011000010000100110 ;
        258:  q   <=  32'b11000000000100001000100011011111 ;
        259:  q   <=  32'b01000000000011101010111100111100 ;
        260:  q   <=  32'b00111110101011001101010100100110 ;
        261:  q   <=  32'b00111111100000000000000111111110 ;
        262:  q   <=  32'b10111111110101010000001101010111 ;
        263:  q   <=  32'b10111111000101110000110010000001 ;
        264:  q   <=  32'b10111110100011100101111001101101 ;
        265:  q   <=  32'b00111110110110000110111000110000 ;
        266:  q   <=  32'b10111111110101011100100100100010 ;
        267:  q   <=  32'b00111110111100010111101000001101 ;
        268:  q   <=  32'b10111111100110110011111010010011 ;
        269:  q   <=  32'b00111101100001111000111010100101 ;
        270:  q   <=  32'b00111111001001110000000011001011 ;
        271:  q   <=  32'b00111110101001110111010001100111 ;
        272:  q   <=  32'b00111111100010101001001110111100 ;
        273:  q   <=  32'b00111111100000001100011100100010 ;
        274:  q   <=  32'b10111111001001101010000111100011 ;
        275:  q   <=  32'b00111110100000111001110011011101 ;
        276:  q   <=  32'b10111111011100011100001010111110 ;
        277:  q   <=  32'b10111111101010010011000001011101 ;
        278:  q   <=  32'b00111111011011001100000101100100 ;
        279:  q   <=  32'b00111000010100010001010100001001 ;
        280:  q   <=  32'b10111101011000001111001010100111 ;
        281:  q   <=  32'b00111111011010010011111110100010 ;
        282:  q   <=  32'b00111111000110000011011010100011 ;
        283:  q   <=  32'b00111110101100110100110110010001 ;
        284:  q   <=  32'b00111111101000000000100000111011 ;
        285:  q   <=  32'b00111111011011100000011010101110 ;
        286:  q   <=  32'b00111110011101011000010001111111 ;
        287:  q   <=  32'b10111111001100001011101110000001 ;
        288:  q   <=  32'b10111111001001101100110000111000 ;
        289:  q   <=  32'b00111111100110001001011011001011 ;
        290:  q   <=  32'b10111111110011100101000001110101 ;
        291:  q   <=  32'b10111100110010000110010001100110 ;
        292:  q   <=  32'b10111111111110010111001111010011 ;
        293:  q   <=  32'b00111111100000101001111110101101 ;
        294:  q   <=  32'b00111111010111001001100101110000 ;
        295:  q   <=  32'b00111010100110000101000100001101 ;
        296:  q   <=  32'b10111101100100010001001100011001 ;
        297:  q   <=  32'b11000000000111110001111101000110 ;
        298:  q   <=  32'b00111111000101001100011110110101 ;
        299:  q   <=  32'b11000000000011000101000011011010 ;
        300:  q   <=  32'b11000000000101000110111100010110 ;
        301:  q   <=  32'b00111101101000111011010001001000 ;
        302:  q   <=  32'b10111111011100101100111110100110 ;
        303:  q   <=  32'b00111110110100101010111011100110 ;
        304:  q   <=  32'b00111111001011010100111001101010 ;
        305:  q   <=  32'b00111111010110111001010001011100 ;
        306:  q   <=  32'b10111111001100001110111111001101 ;
        307:  q   <=  32'b00111110111001100001010011010010 ;
        308:  q   <=  32'b00111101110011100001100011011011 ;
        309:  q   <=  32'b00111111010100110111100101010010 ;
        310:  q   <=  32'b00111111000010010100000110010111 ;
        311:  q   <=  32'b00111111011001011101110000000100 ;
        312:  q   <=  32'b10111110000001110001101010111000 ;
        313:  q   <=  32'b10111110000101101011101111111010 ;
        314:  q   <=  32'b00111111100000001111111010111000 ;
        315:  q   <=  32'b11000000000001111110100111111000 ;
        316:  q   <=  32'b10111111000000010010110010010011 ;
        317:  q   <=  32'b10111111101000101010001011010110 ;
        318:  q   <=  32'b10111110110000111110001000100111 ;
        319:  q   <=  32'b00111111001001100000111111011000 ;
        320:  q   <=  32'b00111111010100110110001011011010 ;
        321:  q   <=  32'b10111111100000011110100110101100 ;
        322:  q   <=  32'b10111110111100010011000000010011 ;
        323:  q   <=  32'b00111110000011000101000000111111 ;
        324:  q   <=  32'b10111110100101010110111100011101 ;
        325:  q   <=  32'b00111110100110101000011111110110 ;
        326:  q   <=  32'b00111110110011001100001110111111 ;
        327:  q   <=  32'b10111111011011100001000111110101 ;
        328:  q   <=  32'b10111110001101010001001011111110 ;
        329:  q   <=  32'b11000000000010000111010000111100 ;
        330:  q   <=  32'b00111111100100101001101100110110 ;
        331:  q   <=  32'b10111111001000010000110000010111 ;
        332:  q   <=  32'b10111111100110100001011111000001 ;
        333:  q   <=  32'b10111110100000100000010100001001 ;
        334:  q   <=  32'b10111111101101101101110111100110 ;
        335:  q   <=  32'b10111100101010101101110110011000 ;
        336:  q   <=  32'b10111111000011111000011110111101 ;
        337:  q   <=  32'b01000000000010110110000010111001 ;
        338:  q   <=  32'b00111111100100011011100100111011 ;
        339:  q   <=  32'b11000000000111111100110011111101 ;
        340:  q   <=  32'b00111110111000011111010110011010 ;
        341:  q   <=  32'b10111111101100101111011000101110 ;
        342:  q   <=  32'b10111110100000101001011010010111 ;
        343:  q   <=  32'b00111110001010000101100110001010 ;
        344:  q   <=  32'b00111111001111110110101101111111 ;
        345:  q   <=  32'b10111110100010111100110011001111 ;
        346:  q   <=  32'b00111111110010011100010000110100 ;
        347:  q   <=  32'b10111110111101100011110101100100 ;
        348:  q   <=  32'b00111110101001111010111110101011 ;
        349:  q   <=  32'b00111111001010100010110000000011 ;
        350:  q   <=  32'b00111101101011100111011101011011 ;
        351:  q   <=  32'b00111111011000011000011000011111 ;
        352:  q   <=  32'b00111110101001010111110000110001 ;
        353:  q   <=  32'b10111111010010001011110111001101 ;
        354:  q   <=  32'b10111111111001110001011001111001 ;
        355:  q   <=  32'b00111111111011011110011001011111 ;
        356:  q   <=  32'b10111111000110101100001001111011 ;
        357:  q   <=  32'b00111101110100111010111001000011 ;
        358:  q   <=  32'b00111111000100000010101110110101 ;
        359:  q   <=  32'b00111101111010001010010110001010 ;
        360:  q   <=  32'b10111111011001111001110000100011 ;
        361:  q   <=  32'b10111110111011110111100001001001 ;
        362:  q   <=  32'b10111101111111111100011001001100 ;
        363:  q   <=  32'b00111111101111010100111010000011 ;
        364:  q   <=  32'b10111111010111000101111001101010 ;
        365:  q   <=  32'b00111111010010001110000000001000 ;
        366:  q   <=  32'b00111110100111100000001111011010 ;
        367:  q   <=  32'b10111110011011110111100100000001 ;
        368:  q   <=  32'b10111111100001110100101011100010 ;
        369:  q   <=  32'b10111110100100010111101011101100 ;
        370:  q   <=  32'b10111101101100011000101010101100 ;
        371:  q   <=  32'b10111111101111000001010100100011 ;
        372:  q   <=  32'b00111110010001001100101101101100 ;
        373:  q   <=  32'b10111111010100101000000111001111 ;
        374:  q   <=  32'b10111101110000010000000100110101 ;
        375:  q   <=  32'b00111110101011000010010000100111 ;
        376:  q   <=  32'b10111111011001111001011101101000 ;
        377:  q   <=  32'b10111110100100111001011001010110 ;
        378:  q   <=  32'b00111110101100110011101101101100 ;
        379:  q   <=  32'b10111111111010101111110101101110 ;
        380:  q   <=  32'b00111111100001001001101011011011 ;
        381:  q   <=  32'b01000000000110110010101001011111 ;
        382:  q   <=  32'b00111111011101011001101101000101 ;
        383:  q   <=  32'b10111110101000011010110011011101 ;
        384:  q   <=  32'b00111110110110110111010001101110 ;
        385:  q   <=  32'b10111111100001001001101100100110 ;
        386:  q   <=  32'b00111111111100000101110111100101 ;
        387:  q   <=  32'b00111111011100001101001000000000 ;
        388:  q   <=  32'b00111111010010011000111101111110 ;
        389:  q   <=  32'b10111111011000000011100101001011 ;
        390:  q   <=  32'b00111110101000111101000001011111 ;
        391:  q   <=  32'b10111111000011101110110001011111 ;
        392:  q   <=  32'b10111110100111110111001110101101 ;
        393:  q   <=  32'b10111111000100011110110000101011 ;
        394:  q   <=  32'b10111111100000110100101100111101 ;
        395:  q   <=  32'b10111111011010001010001110001101 ;
        396:  q   <=  32'b10111110010101101110111101010011 ;
        397:  q   <=  32'b10111111110110010111010001100000 ;
        398:  q   <=  32'b00111111000110111000101110110110 ;
        399:  q   <=  32'b10111101111100010100000000111010 ;
        400:  q   <=  32'b00111111001100101111110000101011 ;
        401:  q   <=  32'b00111110100010100000111101100011 ;
        402:  q   <=  32'b00111110111111010001001100110001 ;
        403:  q   <=  32'b10111111101111011101011011101000 ;
        404:  q   <=  32'b10111111100000101001100000000101 ;
        405:  q   <=  32'b10111110111001001101110010000111 ;
        406:  q   <=  32'b00111101111000001001010010101110 ;
        407:  q   <=  32'b00111111100100000111101001101111 ;
        408:  q   <=  32'b10111110100101000111011000001001 ;
        409:  q   <=  32'b00111111101000010111101001111110 ;
        410:  q   <=  32'b00111110111100110110101011100001 ;
        411:  q   <=  32'b00111111100101100100100101110101 ;
        412:  q   <=  32'b00111110000000011111111001101001 ;
        413:  q   <=  32'b10111111001010000010010100010110 ;
        414:  q   <=  32'b10111111101111011001111001111100 ;
        415:  q   <=  32'b00111110000111110011100010000001 ;
        416:  q   <=  32'b00111111010100011000110010010101 ;
        417:  q   <=  32'b10111110100101011100111000011100 ;
        418:  q   <=  32'b10111111000010100111000011111010 ;
        419:  q   <=  32'b10111110100111100000011001001100 ;
        420:  q   <=  32'b10111111100011000101110100101011 ;
        421:  q   <=  32'b10111110111111000110101111001000 ;
        422:  q   <=  32'b10111110001110010001001110111100 ;
        423:  q   <=  32'b00111101001110111100001111100010 ;
        424:  q   <=  32'b10111101100000101010000010111001 ;
        425:  q   <=  32'b00111111000111001000000001110110 ;
        426:  q   <=  32'b00111101110111111110000111110100 ;
        427:  q   <=  32'b00111111111010000011000110101000 ;
        428:  q   <=  32'b00111110100111111100000110010110 ;
        429:  q   <=  32'b00111111111001101111100110100110 ;
        430:  q   <=  32'b10111111001110010001111001111101 ;
        431:  q   <=  32'b00111111000001101100101111001001 ;
        432:  q   <=  32'b10111110100001010011111110011001 ;
        433:  q   <=  32'b00111111000110011010001011110000 ;
        434:  q   <=  32'b00111111000110000000101111011001 ;
        435:  q   <=  32'b11000000000010111110011111000111 ;
        436:  q   <=  32'b10111111101010011101110010001100 ;
        437:  q   <=  32'b10111111101110000111001100100010 ;
        438:  q   <=  32'b00111110110011011011111010001111 ;
        439:  q   <=  32'b00111111101111000010111110001110 ;
        440:  q   <=  32'b10111110101001110101010000110001 ;
        441:  q   <=  32'b00111111010011111111010001100110 ;
        442:  q   <=  32'b00111111000010111010100010000100 ;
        443:  q   <=  32'b10111111100001101001101111100011 ;
        444:  q   <=  32'b00111110110010111000000011001011 ;
        445:  q   <=  32'b10111111010000000111110000101100 ;
        446:  q   <=  32'b00111111110000100001010100001000 ;
        447:  q   <=  32'b10111101000001010110010001110101 ;
        448:  q   <=  32'b00111111110100010110100001101111 ;
        449:  q   <=  32'b10111110110110011010000101000100 ;
        450:  q   <=  32'b00111111000101101110010100011010 ;
        451:  q   <=  32'b10111101100000001001100010101111 ;
        452:  q   <=  32'b11000000000000010110011111000110 ;
        453:  q   <=  32'b10111111011110110110110011111000 ;
        454:  q   <=  32'b00111111000111001100110110001010 ;
        455:  q   <=  32'b10111101011000001101000001000111 ;
        456:  q   <=  32'b10111111100011110011001010011100 ;
        457:  q   <=  32'b10111111001000000101101001011000 ;
        458:  q   <=  32'b00111110011111111000000110010100 ;
        459:  q   <=  32'b10111111011111100011011001111110 ;
        460:  q   <=  32'b00111111011110011001011001010110 ;
        461:  q   <=  32'b10111111001001000000010110001001 ;
        462:  q   <=  32'b00111111111001111000100011001111 ;
        463:  q   <=  32'b10111111100010100011100100001110 ;
        464:  q   <=  32'b00111110010010111111100001010001 ;
        465:  q   <=  32'b10111111110000101011000011111111 ;
        466:  q   <=  32'b10111111001110010011111111100011 ;
        467:  q   <=  32'b10111111000101111101111101000000 ;
        468:  q   <=  32'b00111110110011010111101111110100 ;
        469:  q   <=  32'b00111111011100010010111110100110 ;
        470:  q   <=  32'b00111110100110011101100101001011 ;
        471:  q   <=  32'b10111110101111110000001100011110 ;
        472:  q   <=  32'b00111111010100001100001111011010 ;
        473:  q   <=  32'b00111111010011001000001111011011 ;
        474:  q   <=  32'b00111101111101100010111000101111 ;
        475:  q   <=  32'b00111111000100100011110101001000 ;
        476:  q   <=  32'b00111110110100110101100111111111 ;
        477:  q   <=  32'b10111111011111001010100110001000 ;
        478:  q   <=  32'b00111111010000100111001100010001 ;
        479:  q   <=  32'b10111111001010000011111001011000 ;
        480:  q   <=  32'b10111111000110101001101001100110 ;
        481:  q   <=  32'b00111110001101010011000110001100 ;
        482:  q   <=  32'b10111110100111010111000100011000 ;
        483:  q   <=  32'b10111110000001101111101111101010 ;
        484:  q   <=  32'b00111111000110000110100101011100 ;
        485:  q   <=  32'b00111111100001011111111010011101 ;
        486:  q   <=  32'b10111110010010101011010110101010 ;
        487:  q   <=  32'b00111110101001111100010101101110 ;
        488:  q   <=  32'b10111110011101000000010101001111 ;
        489:  q   <=  32'b00111110011010110001101101110010 ;
        490:  q   <=  32'b00111110111000010100011101100111 ;
        491:  q   <=  32'b10111111000111011110101011101100 ;
        492:  q   <=  32'b00111110100011001011011101101000 ;
        493:  q   <=  32'b00111111000110011110000111010010 ;
        494:  q   <=  32'b00111101101111010000101111110011 ;
        495:  q   <=  32'b00111111110111010110101101110001 ;
        496:  q   <=  32'b10111111000110111100101001101011 ;
        497:  q   <=  32'b10111111001111001010111111110010 ;
        498:  q   <=  32'b10111111110111111111110000001011 ;
        499:  q   <=  32'b00111111011010010001010101100010 ;
        500:  q   <=  32'b00111111010111011111100100011111 ;
        501:  q   <=  32'b10111101101000111001111011011011 ;
        502:  q   <=  32'b00111111011001100000001010000101 ;
        503:  q   <=  32'b00111110001111000001110011000000 ;
        504:  q   <=  32'b00111110100101001110001001110001 ;
        505:  q   <=  32'b00111101111001110100111110001111 ;
        506:  q   <=  32'b00111110111000010100000101101001 ;
        507:  q   <=  32'b00111101110100000011010001100110 ;
        508:  q   <=  32'b01000000001100100110001110110011 ;
        509:  q   <=  32'b10111111100101010101010101000111 ;
        510:  q   <=  32'b10111111111011010101100110101100 ;
        511:  q   <=  32'b10111111100100100000000111010110 ;
        512:  q   <=  32'b10111111100010111111001010101101 ;
        513:  q   <=  32'b10111110110111100000001000001001 ;
        514:  q   <=  32'b10111110001011001000001101011110 ;
        515:  q   <=  32'b10111110010111111100011101000010 ;
        516:  q   <=  32'b00111111000010101001010011100100 ;
        517:  q   <=  32'b00111110110001110100110111100110 ;
        518:  q   <=  32'b00111111010000000101000010001010 ;
        519:  q   <=  32'b00111111111000111001110111100011 ;
        520:  q   <=  32'b00111111100111001000110101010000 ;
        521:  q   <=  32'b10111111101001000100000110111100 ;
        522:  q   <=  32'b11000000000101010000110110010111 ;
        523:  q   <=  32'b00111111011001101110010011111011 ;
        524:  q   <=  32'b10111111111010101111011000110101 ;
        525:  q   <=  32'b00111101100010001011011111011000 ;
        526:  q   <=  32'b00111101000100010101001011101111 ;
        527:  q   <=  32'b01000000000011101000100111101011 ;
        528:  q   <=  32'b10111101100011011100000000110011 ;
        529:  q   <=  32'b10111111000000011101111111101100 ;
        530:  q   <=  32'b00111110011100010111100000010111 ;
        531:  q   <=  32'b00111110011110111011010001000100 ;
        532:  q   <=  32'b00111101100011110111001111011100 ;
        533:  q   <=  32'b10111111000110111100101111101110 ;
        534:  q   <=  32'b10111111100111000111110111110000 ;
        535:  q   <=  32'b00111110101000100000110001010101 ;
        536:  q   <=  32'b10111111101010111110001100100011 ;
        537:  q   <=  32'b10111111100001000001111010011101 ;
        538:  q   <=  32'b00111111101010100110010101001000 ;
        539:  q   <=  32'b10111110110101100111101001111010 ;
        540:  q   <=  32'b10111110000011111011000001111111 ;
        541:  q   <=  32'b00111111011001100101101011000001 ;
        542:  q   <=  32'b10111110100110011010100000100110 ;
        543:  q   <=  32'b00111111100000111100001001000001 ;
        544:  q   <=  32'b10111110101100001010110001111100 ;
        545:  q   <=  32'b00111111100000011010001101111101 ;
        546:  q   <=  32'b00111111001000010001110000010010 ;
        547:  q   <=  32'b10111110010110100010000010100000 ;
        548:  q   <=  32'b10111111010111011001111001010110 ;
        549:  q   <=  32'b10111111100001011000010010010010 ;
        550:  q   <=  32'b10111110100010100100011001110101 ;
        551:  q   <=  32'b10111110111000000101010000010000 ;
        552:  q   <=  32'b10111110110100010011110111000010 ;
        553:  q   <=  32'b00111111011110111100100110011110 ;
        554:  q   <=  32'b10111110100110000110101111000010 ;
        555:  q   <=  32'b00111111100100100110010000010010 ;
        556:  q   <=  32'b10111111000010000001100001000001 ;
        557:  q   <=  32'b00111111011110001111101000010001 ;
        558:  q   <=  32'b10111111000001011011001000110101 ;
        559:  q   <=  32'b00111110001101001101000011001111 ;
        560:  q   <=  32'b00111111011110001000001001000110 ;
        561:  q   <=  32'b10111110110100111111010000101100 ;
        562:  q   <=  32'b10111110111000000110010011111110 ;
        563:  q   <=  32'b01000000000000000011011110001101 ;
        564:  q   <=  32'b00111111011100110111010001001111 ;
        565:  q   <=  32'b10111110110111010010111110011011 ;
        566:  q   <=  32'b00111111001001100010000011111010 ;
        567:  q   <=  32'b10111110101110000101101111101011 ;
        568:  q   <=  32'b00111111001101001011010011100001 ;
        569:  q   <=  32'b00111111101101010011101010001010 ;
        570:  q   <=  32'b10111111110011010110000011000100 ;
        571:  q   <=  32'b00111111100000111011000101110101 ;
        572:  q   <=  32'b00111111101110101001111010110000 ;
        573:  q   <=  32'b00111101010000100111000101001010 ;
        574:  q   <=  32'b00111111110111111000010101010111 ;
        575:  q   <=  32'b00111110000111110001110111100111 ;
        576:  q   <=  32'b10111111100111100101100111110000 ;
        577:  q   <=  32'b11000000000011000110001000110101 ;
        578:  q   <=  32'b10111110101010101011010001010100 ;
        579:  q   <=  32'b00111111001101101010101011000110 ;
        580:  q   <=  32'b00111110101000101000001101000100 ;
        581:  q   <=  32'b00111110110100111100010010111101 ;
        582:  q   <=  32'b10111111000100111011101111100001 ;
        583:  q   <=  32'b00111110000100110111010100110101 ;
        584:  q   <=  32'b10111111110100011011111111001100 ;
        585:  q   <=  32'b10111111010000101001010101000010 ;
        586:  q   <=  32'b10111111010100011001110001101100 ;
        587:  q   <=  32'b00111111000001010000110011110011 ;
        588:  q   <=  32'b10111100011001111111111110010111 ;
        589:  q   <=  32'b10111111100100111110100001100010 ;
        590:  q   <=  32'b10111100000111000000111001100100 ;
        591:  q   <=  32'b10111111001100001001011101101100 ;
        592:  q   <=  32'b10111111001010101010110011001011 ;
        593:  q   <=  32'b00111111010111010011100011100101 ;
        594:  q   <=  32'b00111101111010000100100001110011 ;
        595:  q   <=  32'b00111110110010111111011000110111 ;
        596:  q   <=  32'b00111111011000100100101111011001 ;
        597:  q   <=  32'b00111110001110001001010101111001 ;
        598:  q   <=  32'b00111111000011010000010011001101 ;
        599:  q   <=  32'b00111111001011101101011010111111 ;
        600:  q   <=  32'b00111111100101011101011010000001 ;
        601:  q   <=  32'b00111110111100111010001111111111 ;
        602:  q   <=  32'b00111111101101001100010000001010 ;
        603:  q   <=  32'b00111100101110010011010101101101 ;
        604:  q   <=  32'b10111101010001000001001010110110 ;
        605:  q   <=  32'b00111111110110011100010101010101 ;
        606:  q   <=  32'b10111111000000100111110001110111 ;
        607:  q   <=  32'b10111011001110110001101001001000 ;
        608:  q   <=  32'b00111111011010110111110001101000 ;
        609:  q   <=  32'b00111110000110010110011101110101 ;
        610:  q   <=  32'b00111111101100111101010011011011 ;
        611:  q   <=  32'b00111111100001000101111000011000 ;
        612:  q   <=  32'b00111110100101010100100010110011 ;
        613:  q   <=  32'b10111111010001110001011101000000 ;
        614:  q   <=  32'b00111111000100010001001011111110 ;
        615:  q   <=  32'b10111111101100001111100110111010 ;
        616:  q   <=  32'b00111110011110100101011110010001 ;
        617:  q   <=  32'b00111111010011101111010111011000 ;
        618:  q   <=  32'b00111110010110100010011110011010 ;
        619:  q   <=  32'b00111111011000010011001010000101 ;
        620:  q   <=  32'b01000000000000100111110011110010 ;
        621:  q   <=  32'b00111111011011001000011011010110 ;
        622:  q   <=  32'b00111110100010001010100101100111 ;
        623:  q   <=  32'b00111111001001000100001111101101 ;
        624:  q   <=  32'b00111110110110011101100100110111 ;
        625:  q   <=  32'b10111111101010000100100011011100 ;
        626:  q   <=  32'b10111110110101010011001111011001 ;
        627:  q   <=  32'b00111111100111001100001010010010 ;
        628:  q   <=  32'b10111101001100101000010101011010 ;
        629:  q   <=  32'b00111111000101010001100110110001 ;
        630:  q   <=  32'b10111111100000001101010011111110 ;
        631:  q   <=  32'b00111101100001000010000101011010 ;
        632:  q   <=  32'b00111111000110011010110010111011 ;
        633:  q   <=  32'b10111111101011100100011000011111 ;
        634:  q   <=  32'b00111110101100011111011110101001 ;
        635:  q   <=  32'b10111110001110100011010100011011 ;
        636:  q   <=  32'b10111111011100001000010101011001 ;
        637:  q   <=  32'b10111101000110011011110001100110 ;
        638:  q   <=  32'b10111111111100101011101000011011 ;
        639:  q   <=  32'b11000000000010000011000011000101 ;
        640:  q   <=  32'b10111111100101101010010101101100 ;
        641:  q   <=  32'b10111111011111011001001110000101 ;
        642:  q   <=  32'b10111111100101100010010111101100 ;
        643:  q   <=  32'b10111111110111001101101011010001 ;
        644:  q   <=  32'b00111110100100111001001010100001 ;
        645:  q   <=  32'b10111111110011000000111000110110 ;
        646:  q   <=  32'b00111101111000011011101001101011 ;
        647:  q   <=  32'b00111111010010010111110100110011 ;
        648:  q   <=  32'b10111011000100011110111101000110 ;
        649:  q   <=  32'b00111101101111101010111111001110 ;
        650:  q   <=  32'b10111110110000011001110111001101 ;
        651:  q   <=  32'b10111111101111011100100001010100 ;
        652:  q   <=  32'b10111101001100110111101100011101 ;
        653:  q   <=  32'b00111111011101011111100010100100 ;
        654:  q   <=  32'b00111111110111100111111011001111 ;
        655:  q   <=  32'b10111110110111000100001111111110 ;
        656:  q   <=  32'b10111111110100000100110000011100 ;
        657:  q   <=  32'b00111110001010100101011011111111 ;
        658:  q   <=  32'b00111110110000001010010111101100 ;
        659:  q   <=  32'b10111110011010000110010110110011 ;
        660:  q   <=  32'b10111111100100110000111110001110 ;
        661:  q   <=  32'b01000000000000011000111010101010 ;
        662:  q   <=  32'b11000000000101110000001001101110 ;
        663:  q   <=  32'b10111111000000101000110110000111 ;
        664:  q   <=  32'b10111111101010010010101100000111 ;
        665:  q   <=  32'b10111111001000101101100101001101 ;
        666:  q   <=  32'b00111110101000101011110101101011 ;
        667:  q   <=  32'b00111110000011010101110001110010 ;
        668:  q   <=  32'b10111111001101011111001010111011 ;
        669:  q   <=  32'b00111111010001101110100110110100 ;
        670:  q   <=  32'b00111111000111110101010100110101 ;
        671:  q   <=  32'b00111111001001011011101011000000 ;
        672:  q   <=  32'b10111110110110011110110001100101 ;
        673:  q   <=  32'b00111111100001100011011111100100 ;
        674:  q   <=  32'b00111111001010010010010000011001 ;
        675:  q   <=  32'b01000000001000001000111110111010 ;
        676:  q   <=  32'b00111111100010000001111101110010 ;
        677:  q   <=  32'b00111111100101000001011000000010 ;
        678:  q   <=  32'b00111101010110010000000001010011 ;
        679:  q   <=  32'b10111111101001001110100111010101 ;
        680:  q   <=  32'b10111110101111100001000010110110 ;
        681:  q   <=  32'b10111111010000011111111010100110 ;
        682:  q   <=  32'b10111111000100000110000001000100 ;
        683:  q   <=  32'b00111111000011100001110110001111 ;
        684:  q   <=  32'b10111111000011101000100100000001 ;
        685:  q   <=  32'b10111111011001010010011000100010 ;
        686:  q   <=  32'b10111110110100011001001101100111 ;
        687:  q   <=  32'b10111110001001001011111110000000 ;
        688:  q   <=  32'b00111110110100011001010001001000 ;
        689:  q   <=  32'b10111111011100111101111111110011 ;
        690:  q   <=  32'b00111110101000100111011101101111 ;
        691:  q   <=  32'b00111101100111111100100011111110 ;
        692:  q   <=  32'b00111111101010011000010101110110 ;
        693:  q   <=  32'b10111110010110100100100101011101 ;
        694:  q   <=  32'b10111110000010011011010011000101 ;
        695:  q   <=  32'b10111111100101011110111011111100 ;
        696:  q   <=  32'b10111111101100010101000001001001 ;
        697:  q   <=  32'b00111110100111101111101011110010 ;
        698:  q   <=  32'b10111110011111110111101000001111 ;
        699:  q   <=  32'b00111111000000001111010101011110 ;
        700:  q   <=  32'b10111111011001001000010101110101 ;
        701:  q   <=  32'b00111111111101000100101000100001 ;
        702:  q   <=  32'b00111101111110100101010000010110 ;
        703:  q   <=  32'b00111111100001100000010100101111 ;
        704:  q   <=  32'b10111110011010000101110111000100 ;
        705:  q   <=  32'b10111110001001100110011011101000 ;
        706:  q   <=  32'b00111111001100001010011100111101 ;
        707:  q   <=  32'b00111111000011100100011000010011 ;
        708:  q   <=  32'b10111111100011110110010010000100 ;
        709:  q   <=  32'b10111111110001000010111101001000 ;
        710:  q   <=  32'b10111111100011001000011011101110 ;
        711:  q   <=  32'b10111111101101010011100000001111 ;
        712:  q   <=  32'b00111101011101000000000001001010 ;
        713:  q   <=  32'b10111110110100101000111101111011 ;
        714:  q   <=  32'b10111110101111000110101111100111 ;
        715:  q   <=  32'b10111111101011100011010000001010 ;
        716:  q   <=  32'b00111111010001111001000110111011 ;
        717:  q   <=  32'b00111110111000001111101001111110 ;
        718:  q   <=  32'b10111101101101111000101111111110 ;
        719:  q   <=  32'b00111111100000101011011000000111 ;
        720:  q   <=  32'b10111111010111111011110100011110 ;
        721:  q   <=  32'b00111110110101000101001110011000 ;
        722:  q   <=  32'b00111110101100100110011011100010 ;
        723:  q   <=  32'b00111110101100101101000101111001 ;
        724:  q   <=  32'b10111111001110101010111111110010 ;
        725:  q   <=  32'b00111110101001110101011110011010 ;
        726:  q   <=  32'b10111111000000111100111101001000 ;
        727:  q   <=  32'b10111111011001010111110101111110 ;
        728:  q   <=  32'b10111111100110100000010010110001 ;
        729:  q   <=  32'b00111111100001001101011100100100 ;
        730:  q   <=  32'b10111111010110001000111111001100 ;
        731:  q   <=  32'b10111110001100010001000001010011 ;
        732:  q   <=  32'b10111111100110101011010100011100 ;
        733:  q   <=  32'b10111110100110000010000100000001 ;
        734:  q   <=  32'b11000000010011101101100110110101 ;
        735:  q   <=  32'b10111111100010110010000101111010 ;
        736:  q   <=  32'b10111111101101101001010101110101 ;
        737:  q   <=  32'b10111111100000011101100110000101 ;
        738:  q   <=  32'b10111110010110100110001010110110 ;
        739:  q   <=  32'b10111110101001101001001111111011 ;
        740:  q   <=  32'b00111111111110001110001000000110 ;
        741:  q   <=  32'b10111111000100100101111110111010 ;
        742:  q   <=  32'b10111110100000000000010000111011 ;
        743:  q   <=  32'b10111111110010001101111101010100 ;
        744:  q   <=  32'b10111110111101000110101110000000 ;
        745:  q   <=  32'b10111111101010110100001011010001 ;
        746:  q   <=  32'b00111100111110000011010110101000 ;
        747:  q   <=  32'b00111111010110100110001111100100 ;
        748:  q   <=  32'b00111110110011101111101001001111 ;
        749:  q   <=  32'b10111111001100110101101111011000 ;
        750:  q   <=  32'b10111111110100001011010110100001 ;
        751:  q   <=  32'b00111111101110101110000110110110 ;
        752:  q   <=  32'b01000000000000110011001111100110 ;
        753:  q   <=  32'b00111101111101101100100100000100 ;
        754:  q   <=  32'b10111111011111010110101000110001 ;
        755:  q   <=  32'b00111111100110010101000010010011 ;
        756:  q   <=  32'b10111111000101111011100001010001 ;
        757:  q   <=  32'b10111110111100001000101011011010 ;
        758:  q   <=  32'b00111111011000101110100110100000 ;
        759:  q   <=  32'b10111111101100010100111011100001 ;
        760:  q   <=  32'b10111111111110100111011011101001 ;
        761:  q   <=  32'b00111110110101110110001111011010 ;
        762:  q   <=  32'b00111110110011010010110110000111 ;
        763:  q   <=  32'b00111101110000101101100111100100 ;
        764:  q   <=  32'b00111110111111100100110101101010 ;
        765:  q   <=  32'b00111111100010101000011011011100 ;
        766:  q   <=  32'b00111111011110000110111101000100 ;
        767:  q   <=  32'b10111111000100011000110111000110 ;
        768:  q   <=  32'b00111111010011110101101001010100 ;
        769:  q   <=  32'b00111110001100010110011111000010 ;
        770:  q   <=  32'b10111111000000010110101100111100 ;
        771:  q   <=  32'b10111111100110001011111000111110 ;
        772:  q   <=  32'b00111111001001011001111111100011 ;
        773:  q   <=  32'b10111110101101010000111000000101 ;
        774:  q   <=  32'b00111101001111100011001000100001 ;
        775:  q   <=  32'b10111111010010101111111010011011 ;
        776:  q   <=  32'b10111111110001100111011101000010 ;
        777:  q   <=  32'b00111110001011111011010001010101 ;
        778:  q   <=  32'b10111101011111101000010110011000 ;
        779:  q   <=  32'b00111111100110010111100110111110 ;
        780:  q   <=  32'b00111111010011010011110001111010 ;
        781:  q   <=  32'b00111111100001101101001010101111 ;
        782:  q   <=  32'b10111111001111111011011001100011 ;
        783:  q   <=  32'b10111111011011111011001100010111 ;
        784:  q   <=  32'b10111111101000100111000101101111 ;
        785:  q   <=  32'b00111110111111101111011101010000 ;
        786:  q   <=  32'b01000000001100101000000001001110 ;
        787:  q   <=  32'b00111111001110100100001000101001 ;
        788:  q   <=  32'b10111111010001011110011110000111 ;
        789:  q   <=  32'b00111111010101100010110110100001 ;
        790:  q   <=  32'b10111111100100000110110100100000 ;
        791:  q   <=  32'b10111111101101100101010100001001 ;
        792:  q   <=  32'b00111111001101111010101001001100 ;
        793:  q   <=  32'b10111111010001110010010011010000 ;
        794:  q   <=  32'b00111110101000011100100011100110 ;
        795:  q   <=  32'b00111111101101000000100101010111 ;
        796:  q   <=  32'b00111110110011010110000000110101 ;
        797:  q   <=  32'b00111111011011011111111000110111 ;
        798:  q   <=  32'b10111111110011011000101011101101 ;
        799:  q   <=  32'b00111111001010010101101001110000 ;
        800:  q   <=  32'b01000000000010001101110100111000 ;
        801:  q   <=  32'b00111111000010101000100000011100 ;
        802:  q   <=  32'b10111111110001010011101101110110 ;
        803:  q   <=  32'b10111110010100000000010010101010 ;
        804:  q   <=  32'b10111110111111111111101101110001 ;
        805:  q   <=  32'b00111110110001000001101110110101 ;
        806:  q   <=  32'b00111110110100101111011001001101 ;
        807:  q   <=  32'b00111110110011111001110010111000 ;
        808:  q   <=  32'b10111110101110100100000101111000 ;
        809:  q   <=  32'b10111111000110010110100111100100 ;
        810:  q   <=  32'b10111111000101101110111101001101 ;
        811:  q   <=  32'b00111111010110101000000110100110 ;
        812:  q   <=  32'b10111111111011010010111101011110 ;
        813:  q   <=  32'b10111110010101000100011101000111 ;
        814:  q   <=  32'b00111110100010100110111100000011 ;
        815:  q   <=  32'b10111111001001110001110000000000 ;
        816:  q   <=  32'b00111110111101000101011100100010 ;
        817:  q   <=  32'b10111101100100100001000000001001 ;
        818:  q   <=  32'b10111111011100000011010010000011 ;
        819:  q   <=  32'b00111110001001010011110001111011 ;
        820:  q   <=  32'b10111110100010010100111101000100 ;
        821:  q   <=  32'b10111110110100011101101011010011 ;
        822:  q   <=  32'b10111111001101100001100100111110 ;
        823:  q   <=  32'b00111101011110111010111001000010 ;
        824:  q   <=  32'b10111111111011000100110111110110 ;
        825:  q   <=  32'b10111110110010111111001001010001 ;
        826:  q   <=  32'b10111111000010110010010111111000 ;
        827:  q   <=  32'b10111111011010010111001000101110 ;
        828:  q   <=  32'b00111111001001110001011101000001 ;
        829:  q   <=  32'b10111111001110111111100100110011 ;
        830:  q   <=  32'b00111111000010100110011011101110 ;
        831:  q   <=  32'b00111111011110011101000010110101 ;
        832:  q   <=  32'b10111110001000001010001010100011 ;
        833:  q   <=  32'b00111110100011100011101110110110 ;
        834:  q   <=  32'b00111111001000111011011101100111 ;
        835:  q   <=  32'b10111101101001011101011111001101 ;
        836:  q   <=  32'b00111111000010100111011001110111 ;
        837:  q   <=  32'b10111111101000011001101110111001 ;
        838:  q   <=  32'b00111111100011100010001001011110 ;
        839:  q   <=  32'b10111111011111010101001111111010 ;
        840:  q   <=  32'b10111111111010100001011101001011 ;
        841:  q   <=  32'b00111111101100010011011100111111 ;
        842:  q   <=  32'b10111101100000000111011011100111 ;
        843:  q   <=  32'b00111110111001011101100011111101 ;
        844:  q   <=  32'b10111110101110011111110100000011 ;
        845:  q   <=  32'b10111111100000101010001001111010 ;
        846:  q   <=  32'b11000000010001001010101111011000 ;
        847:  q   <=  32'b00111111001000000101001111010010 ;
        848:  q   <=  32'b10111110100100101100100001010000 ;
        849:  q   <=  32'b10111110010010100001010001000010 ;
        850:  q   <=  32'b00111110110011111010101110000001 ;
        851:  q   <=  32'b10111111101101011010110100110101 ;
        852:  q   <=  32'b10111111001110101011110011101100 ;
        853:  q   <=  32'b00111111100100101101101110100011 ;
        854:  q   <=  32'b00111111000110010000110110101000 ;
        855:  q   <=  32'b10111111101001000000000100000110 ;
        856:  q   <=  32'b11000000000011010000001001001000 ;
        857:  q   <=  32'b10111111000100100011110100110010 ;
        858:  q   <=  32'b00111110010110110010000111100100 ;
        859:  q   <=  32'b00111111011100010011111110011101 ;
        860:  q   <=  32'b00111101101111111111001100100110 ;
        861:  q   <=  32'b10111111100011111010011111101001 ;
        862:  q   <=  32'b00111110100111001100000010110111 ;
        863:  q   <=  32'b10111111100101100000111100010001 ;
        864:  q   <=  32'b10111111011101100000000111100111 ;
        865:  q   <=  32'b10111111001001110101101100101101 ;
        866:  q   <=  32'b10111111100111010101110011000101 ;
        867:  q   <=  32'b10111110100010101011101111110001 ;
        868:  q   <=  32'b10111111011001100110001100100000 ;
        869:  q   <=  32'b10111110100100100100010101110100 ;
        870:  q   <=  32'b10111110111011001100001010000100 ;
        871:  q   <=  32'b10111110110100011100111101011110 ;
        872:  q   <=  32'b10111111000000001110011111101110 ;
        873:  q   <=  32'b00111111100111011101110010101110 ;
        874:  q   <=  32'b00111111000111000011110011110110 ;
        875:  q   <=  32'b00111101011100011111010110100100 ;
        876:  q   <=  32'b10111111101110111100010011101001 ;
        877:  q   <=  32'b10111111110100000001101001010010 ;
        878:  q   <=  32'b10111111111110110111110100000001 ;
        879:  q   <=  32'b01000000001001101011101110000110 ;
        880:  q   <=  32'b00111111011110001110110110001110 ;
        881:  q   <=  32'b00111110100000111001001100000010 ;
        882:  q   <=  32'b10111111011110010110011111010010 ;
        883:  q   <=  32'b10111111100100101011110000010001 ;
        884:  q   <=  32'b00111111000011000011001000011010 ;
        885:  q   <=  32'b00111111110010000101010010101100 ;
        886:  q   <=  32'b10111111110110001011111101111100 ;
        887:  q   <=  32'b10111110111001100001011101101001 ;
        888:  q   <=  32'b10111101101011001010000101010010 ;
        889:  q   <=  32'b10111111111111101111100111000011 ;
        890:  q   <=  32'b00111111010101110101101111100000 ;
        891:  q   <=  32'b10111110110101000100111000101100 ;
        892:  q   <=  32'b00111111111101001100001001010111 ;
        893:  q   <=  32'b10111110110010000010001111100000 ;
        894:  q   <=  32'b00111110110100011000000001010000 ;
        895:  q   <=  32'b10111111100100100011101100010110 ;
        896:  q   <=  32'b10111111000111111111011100010010 ;
        897:  q   <=  32'b10111111100101011001100010110101 ;
        898:  q   <=  32'b00111110110010001111111110100000 ;
        899:  q   <=  32'b00111111101001101010001010101101 ;
        900:  q   <=  32'b10111111000101111111100011101000 ;
        901:  q   <=  32'b00111110110111110110110010011000 ;
        902:  q   <=  32'b10111111000000010001110111100110 ;
        903:  q   <=  32'b00111101110100010001110111011001 ;
        904:  q   <=  32'b00111111100110010001111010111100 ;
        905:  q   <=  32'b00111101111101100101011011010110 ;
        906:  q   <=  32'b10111111100001001011011101001000 ;
        907:  q   <=  32'b10111111010110110110101100011110 ;
        908:  q   <=  32'b10111110001011011111001110000111 ;
        909:  q   <=  32'b10111110010001000100010010110000 ;
        910:  q   <=  32'b10111111010111011010011000010000 ;
        911:  q   <=  32'b00111110001110010000000000000100 ;
        912:  q   <=  32'b00111111101000100001110110011010 ;
        913:  q   <=  32'b10111110100000001001100101000010 ;
        914:  q   <=  32'b10111110010100010111101011001111 ;
        915:  q   <=  32'b11000000000011001110010110111100 ;
        916:  q   <=  32'b10111111010001100100011001111101 ;
        917:  q   <=  32'b10111111101100100101011011000001 ;
        918:  q   <=  32'b10111110110001011100000010001100 ;
        919:  q   <=  32'b00111111000001101000110011010011 ;
        920:  q   <=  32'b00111111110000101111101001111100 ;
        921:  q   <=  32'b00111111111001100011010100010000 ;
        922:  q   <=  32'b10111101111011110110000100000100 ;
        923:  q   <=  32'b10111110101000111111000011000001 ;
        924:  q   <=  32'b00111111010100010100100010111111 ;
        925:  q   <=  32'b00111110111110101111011000100101 ;
        926:  q   <=  32'b00111111010000111110011110000000 ;
        927:  q   <=  32'b00111111010001110011110101001011 ;
        928:  q   <=  32'b10111111101111010111101010100011 ;
        929:  q   <=  32'b00111111000010100101010101001010 ;
        930:  q   <=  32'b10111101101110110111100011001111 ;
        931:  q   <=  32'b10111111010000101001111111100110 ;
        932:  q   <=  32'b10111111001100011000111101111000 ;
        933:  q   <=  32'b00111111101001000000011011001110 ;
        934:  q   <=  32'b10111111010011110100101011110110 ;
        935:  q   <=  32'b10111111100111100101000000010000 ;
        936:  q   <=  32'b00111110010110111101011011000011 ;
        937:  q   <=  32'b01000000000000001011000001111100 ;
        938:  q   <=  32'b00111100110100010101011110000111 ;
        939:  q   <=  32'b00111110100111011101100101101100 ;
        940:  q   <=  32'b10111111011100000011000011111000 ;
        941:  q   <=  32'b00111111110101100100110010110101 ;
        942:  q   <=  32'b00111101111111111111100111001100 ;
        943:  q   <=  32'b00111111000001111011010010110111 ;
        944:  q   <=  32'b10111111011100111011101010111110 ;
        945:  q   <=  32'b00111111010110101010001010001100 ;
        946:  q   <=  32'b00111110110001110011111000011100 ;
        947:  q   <=  32'b10111111100100111111011111010111 ;
        948:  q   <=  32'b00111101001000101100011010001011 ;
        949:  q   <=  32'b10111110111001101011010011011100 ;
        950:  q   <=  32'b00111101110111111011110101100010 ;
        951:  q   <=  32'b10111110100000000100100001110110 ;
        952:  q   <=  32'b10111110010000100111010110010100 ;
        953:  q   <=  32'b10111111100001000011011010000010 ;
        954:  q   <=  32'b10111110101001011000011010000100 ;
        955:  q   <=  32'b00111111010001000011101100011010 ;
        956:  q   <=  32'b00111111110111110101000101110011 ;
        957:  q   <=  32'b10111111100101001000101111101010 ;
        958:  q   <=  32'b01000000000110000010011110000100 ;
        959:  q   <=  32'b00111111110000110101011010000101 ;
        960:  q   <=  32'b00111110001011001000110100111010 ;
        961:  q   <=  32'b10111110100110100011011110111110 ;
        962:  q   <=  32'b10111111001100101101101100000001 ;
        963:  q   <=  32'b00111111010101010011000001110011 ;
        964:  q   <=  32'b10111111001100011101000110100110 ;
        965:  q   <=  32'b10111110111011000111101111101101 ;
        966:  q   <=  32'b00111111011000100011010010111011 ;
        967:  q   <=  32'b00111110110111110011010000010011 ;
        968:  q   <=  32'b00111111011001011001000100111100 ;
        969:  q   <=  32'b00111111000000010011011000011110 ;
        970:  q   <=  32'b10111110110011010100001001100011 ;
        971:  q   <=  32'b10111111000000111000101110001011 ;
        972:  q   <=  32'b00111111010010111101111010111111 ;
        973:  q   <=  32'b10111111001010111101001100011110 ;
        974:  q   <=  32'b00111111100101111110010001110001 ;
        975:  q   <=  32'b00111111010010100110101101110001 ;
        976:  q   <=  32'b00111110100100110101000000111011 ;
        977:  q   <=  32'b00111011010100110110110100111000 ;
        978:  q   <=  32'b00111110101110110011001000101101 ;
        979:  q   <=  32'b01000000011000011011010100010110 ;
        980:  q   <=  32'b10111101111001100100010100110001 ;
        981:  q   <=  32'b10111111110001110011111001111000 ;
        982:  q   <=  32'b00111111111101010010001000010010 ;
        983:  q   <=  32'b00111111000111000001111011011110 ;
        984:  q   <=  32'b10111111001001011101110110001001 ;
        985:  q   <=  32'b01000000001001111000001001101010 ;
        986:  q   <=  32'b00111111000011010000101100010110 ;
        987:  q   <=  32'b00111110100101101010000111011101 ;
        988:  q   <=  32'b10111111010001110010000011000101 ;
        989:  q   <=  32'b10111111100010000100111110100001 ;
        990:  q   <=  32'b10111111111000100101101101100100 ;
        991:  q   <=  32'b10111110110110001000100011101000 ;
        992:  q   <=  32'b10111111100001101100110000001111 ;
        993:  q   <=  32'b00111111001001011101001101001001 ;
        994:  q   <=  32'b10111110101000101010000000101001 ;
        995:  q   <=  32'b00111111111000100110111001010000 ;
        996:  q   <=  32'b00111111110000010101101011000011 ;
        997:  q   <=  32'b00111110001001111111001001010010 ;
        998:  q   <=  32'b10111110100100001100011001100111 ;
        999:  q   <=  32'b00111111100100110111101000101011 ;
        1000:  q   <=  32'b10111111100100101100000011000011 ;
        1001:  q   <=  32'b00111111001011000111011110000100 ;
        1002:  q   <=  32'b10111111001010110100101011111101 ;
        1003:  q   <=  32'b10111110110011001111011100011000 ;
        1004:  q   <=  32'b10111111001010111111101100111110 ;
        1005:  q   <=  32'b00111111000100110101110001101100 ;
        1006:  q   <=  32'b10111111010001110011000100100010 ;
        1007:  q   <=  32'b10111111100010000010001011000110 ;
        1008:  q   <=  32'b00111111000011011000111111111100 ;
        1009:  q   <=  32'b10111110110110001100101110101010 ;
        1010:  q   <=  32'b00111110101110010010000111110011 ;
        1011:  q   <=  32'b10111110101101000010101011010011 ;
        1012:  q   <=  32'b00111110100010100000000100111101 ;
        1013:  q   <=  32'b11000000001001000001111111110000 ;
        1014:  q   <=  32'b00111110111011101000010110111110 ;
        1015:  q   <=  32'b00111111111011010100000101111100 ;
        1016:  q   <=  32'b00111111100001010000011101101110 ;
        1017:  q   <=  32'b00111111011010010011000010000100 ;
        1018:  q   <=  32'b10111110011101010111110000011110 ;
        1019:  q   <=  32'b00111110001110010101011110001111 ;
        1020:  q   <=  32'b00111110011110100001110010001101 ;
        1021:  q   <=  32'b00111101110001010110100110100001 ;
        1022:  q   <=  32'b10111111010101001001100110010101 ;
        1023:  q   <=  32'b10111110101101000101101001100110 ;
        1024:  q   <=  32'b10111110001100101111100000111010 ;
        1025:  q   <=  32'b10111110111101100001100000110100 ;
        1026:  q   <=  32'b00111111010101100011101011101110 ;
        1027:  q   <=  32'b01000000001000100111010001010000 ;
        1028:  q   <=  32'b10111111101010010110001100000100 ;
        1029:  q   <=  32'b00111110000000110110101110100001 ;
        1030:  q   <=  32'b10111111101110001001111111100001 ;
        1031:  q   <=  32'b00111111101001101011100010010110 ;
        1032:  q   <=  32'b00111111101101000111011111111010 ;
        1033:  q   <=  32'b10111111110101001100111000110101 ;
        1034:  q   <=  32'b00111111111110001100101010100111 ;
        1035:  q   <=  32'b10111111100010101101011101100110 ;
        1036:  q   <=  32'b00111110011010000100001100111011 ;
        1037:  q   <=  32'b00111111100011001010100110110110 ;
        1038:  q   <=  32'b00111110000101101011100010100101 ;
        1039:  q   <=  32'b01000000000100101110110000110000 ;
        1040:  q   <=  32'b01000000001100000010100111101000 ;
        1041:  q   <=  32'b00111110000011011010001100101001 ;
        1042:  q   <=  32'b10111111111101000001101010111110 ;
        1043:  q   <=  32'b10111110101110101110000001011100 ;
        1044:  q   <=  32'b10111111010110010001110110111100 ;
        1045:  q   <=  32'b10111111010000111100011011100000 ;
        1046:  q   <=  32'b10111111100100000101100001001101 ;
        1047:  q   <=  32'b00111101101000000010000101111111 ;
        1048:  q   <=  32'b01000000000001101101001100000101 ;
        1049:  q   <=  32'b10111111001101110100000111000110 ;
        1050:  q   <=  32'b10111110100011111001111110111111 ;
        1051:  q   <=  32'b00111111100101010100111100001101 ;
        1052:  q   <=  32'b00111111100110110011110110111011 ;
        1053:  q   <=  32'b00111110111110001001100011010100 ;
        1054:  q   <=  32'b00111111100000110101010010000010 ;
        1055:  q   <=  32'b00111111010111101110011111100110 ;
        1056:  q   <=  32'b10111110110000110111010111000100 ;
        1057:  q   <=  32'b00111110110110111001011111011101 ;
        1058:  q   <=  32'b10111110100110010010011110100010 ;
        1059:  q   <=  32'b10111111011001100101110111001000 ;
        1060:  q   <=  32'b00111111001000100111111010101101 ;
        1061:  q   <=  32'b00111101100010100010010100011011 ;
        1062:  q   <=  32'b10111110001111111001110010000111 ;
        1063:  q   <=  32'b00111110100101010101110101001101 ;
        1064:  q   <=  32'b00111111011111001101100110001111 ;
        1065:  q   <=  32'b00111110110010010010111010111000 ;
        1066:  q   <=  32'b00111110010001110011100001111001 ;
        1067:  q   <=  32'b00111110100011110011111111111001 ;
        1068:  q   <=  32'b00111101010100011100110001100011 ;
        1069:  q   <=  32'b10111111010001100100001101101011 ;
        1070:  q   <=  32'b00111111010010010110101010000110 ;
        1071:  q   <=  32'b00111111101101000101011100010000 ;
        1072:  q   <=  32'b10111111000010001011101010101111 ;
        1073:  q   <=  32'b00111111111101101100000011001001 ;
        1074:  q   <=  32'b10111110001101000111101000111100 ;
        1075:  q   <=  32'b10111110011110011001100110110001 ;
        1076:  q   <=  32'b10111111011001011100100100101000 ;
        1077:  q   <=  32'b10111111010010101101011010010110 ;
        1078:  q   <=  32'b10111111011100111111011000100110 ;
        1079:  q   <=  32'b00111110101101010011001100011000 ;
        1080:  q   <=  32'b00111111110011000110101101011011 ;
        1081:  q   <=  32'b00111111000001110000100001001010 ;
        1082:  q   <=  32'b00111111010110101010110100000000 ;
        1083:  q   <=  32'b00111111101010111100000110100000 ;
        1084:  q   <=  32'b11000000000111111111100001011011 ;
        1085:  q   <=  32'b10111110001010111001010010101011 ;
        1086:  q   <=  32'b00111110101101001011111001101100 ;
        1087:  q   <=  32'b00111111001101111001110111110000 ;
        1088:  q   <=  32'b10111111101001110000010101100000 ;
        1089:  q   <=  32'b10111111100000001100000001010000 ;
        1090:  q   <=  32'b00111111010010100110101000111011 ;
        1091:  q   <=  32'b10111101111011101011110011110010 ;
        1092:  q   <=  32'b00111111000011011001011101001100 ;
        1093:  q   <=  32'b10111111011101011110110011010001 ;
        1094:  q   <=  32'b10111111110100010010000001101111 ;
        1095:  q   <=  32'b00111111010000101101111000000101 ;
        1096:  q   <=  32'b00111111100110001011111001001001 ;
        1097:  q   <=  32'b00111111110100001110011101000000 ;
        1098:  q   <=  32'b10111111110001000001111011001001 ;
        1099:  q   <=  32'b10111111101010110001110111111010 ;
        1100:  q   <=  32'b10111111101111001010011100000000 ;
        1101:  q   <=  32'b10111101001010101010011011100110 ;
        1102:  q   <=  32'b10111111000111011001000111100011 ;
        1103:  q   <=  32'b00111111101010000011011000111001 ;
        1104:  q   <=  32'b10111111101110100011111110011111 ;
        1105:  q   <=  32'b10111111110111110000010101001100 ;
        1106:  q   <=  32'b00111110010100100011101101100100 ;
        1107:  q   <=  32'b00111111100110001011000111110001 ;
        1108:  q   <=  32'b10111111010011011000010111010000 ;
        1109:  q   <=  32'b10111111101000100000000001011111 ;
        1110:  q   <=  32'b10111110000110001110101001010001 ;
        1111:  q   <=  32'b10111111110100010111011100010101 ;
        1112:  q   <=  32'b00111100100011100001010110111010 ;
        1113:  q   <=  32'b00111111010101000001000100110000 ;
        1114:  q   <=  32'b00111110010111101111011011001101 ;
        1115:  q   <=  32'b10111111111101000110001000100011 ;
        1116:  q   <=  32'b10111111000010010110110100100111 ;
        1117:  q   <=  32'b10111110100110101010001111111010 ;
        1118:  q   <=  32'b00111111111010000010001101110101 ;
        1119:  q   <=  32'b00111111011010100011001110111001 ;
        1120:  q   <=  32'b10111101011010011100110101111000 ;
        1121:  q   <=  32'b00111111101001111001100100101101 ;
        1122:  q   <=  32'b10111111100001011011100111100111 ;
        1123:  q   <=  32'b10111110101100100101000000000111 ;
        1124:  q   <=  32'b00111111101101001100111011001101 ;
        1125:  q   <=  32'b00111111110000000100111000010101 ;
        1126:  q   <=  32'b00111111001110101111100111101011 ;
        1127:  q   <=  32'b00111110111110110100001111100001 ;
        1128:  q   <=  32'b10111111000101100000110001011100 ;
        1129:  q   <=  32'b00111111001111101011000110111110 ;
        1130:  q   <=  32'b10111111010101000000000111110110 ;
        1131:  q   <=  32'b00111111000100110001001111001010 ;
        1132:  q   <=  32'b00111110100100000100110110000011 ;
        1133:  q   <=  32'b00111111100100011101010011001001 ;
        1134:  q   <=  32'b10111110110110100000101101011001 ;
        1135:  q   <=  32'b00111111001000101101101000010000 ;
        1136:  q   <=  32'b00111111010010110000110110110111 ;
        1137:  q   <=  32'b10111111011001011111110000001010 ;
        1138:  q   <=  32'b00111110000111111111111010100110 ;
        1139:  q   <=  32'b00111111110011000111001011010000 ;
        1140:  q   <=  32'b00111101111001100100011011001010 ;
        1141:  q   <=  32'b10111110100111100000010000010110 ;
        1142:  q   <=  32'b00111110111010011100111101001001 ;
        1143:  q   <=  32'b10111110100011001101101000000100 ;
        1144:  q   <=  32'b00111110111000101110001110111000 ;
        1145:  q   <=  32'b10111110000010011111111111011110 ;
        1146:  q   <=  32'b10111100100101100010010100010101 ;
        1147:  q   <=  32'b00111110111010111110110010010111 ;
        1148:  q   <=  32'b00111111101011100110000001011010 ;
        1149:  q   <=  32'b00111110111001110101110000011010 ;
        1150:  q   <=  32'b00111111110100101111111000111100 ;
        1151:  q   <=  32'b11000000000000011101000010101110 ;
        1152:  q   <=  32'b10111110111001100000010011111101 ;
        1153:  q   <=  32'b00111110011100011010100000110011 ;
        1154:  q   <=  32'b10111111010101011100110111100101 ;
        1155:  q   <=  32'b10111111101000110101001001111111 ;
        1156:  q   <=  32'b00111111000111011111011000000010 ;
        1157:  q   <=  32'b00111111000111001101101000000001 ;
        1158:  q   <=  32'b00111110100101000010100111000100 ;
        1159:  q   <=  32'b00111110110010100110011011011111 ;
        1160:  q   <=  32'b10111111010111101101110100110100 ;
        1161:  q   <=  32'b10111110111111101101000100000010 ;
        1162:  q   <=  32'b10111101110110100111011011000000 ;
        1163:  q   <=  32'b10111111001100000001010110010001 ;
        1164:  q   <=  32'b00111110101010011110110001001010 ;
        1165:  q   <=  32'b01000000000101110101111111010111 ;
        1166:  q   <=  32'b10111110111101101110011011110001 ;
        1167:  q   <=  32'b00111111001001011011111100101010 ;
        1168:  q   <=  32'b10111111100001000110100000000111 ;
        1169:  q   <=  32'b00111111101010110111011010000110 ;
        1170:  q   <=  32'b10111111011110000001100110010101 ;
        1171:  q   <=  32'b00111110010101011011100110001010 ;
        1172:  q   <=  32'b10111111000111100101110000100010 ;
        1173:  q   <=  32'b00111111000000110001001101110101 ;
        1174:  q   <=  32'b00111100001110100000011011011000 ;
        1175:  q   <=  32'b10111101001101000010110101101010 ;
        1176:  q   <=  32'b01000000001111001011110111101110 ;
        1177:  q   <=  32'b10111111001000010100101010110101 ;
        1178:  q   <=  32'b10111101010000000000010010011100 ;
        1179:  q   <=  32'b01000000001010111011011010110000 ;
        1180:  q   <=  32'b10111111100100101100011011000010 ;
        1181:  q   <=  32'b00111111000011011001000101010011 ;
        1182:  q   <=  32'b10111111100010011100100101100011 ;
        1183:  q   <=  32'b00111111100000111110101111111111 ;
        1184:  q   <=  32'b00111110101001111011000111111100 ;
        1185:  q   <=  32'b00111111001001101111000110100110 ;
        1186:  q   <=  32'b10111110100011101100011011100010 ;
        1187:  q   <=  32'b00111110011110110001001110000001 ;
        1188:  q   <=  32'b00111111101111000111101101010010 ;
        1189:  q   <=  32'b11000000000100011001101101000011 ;
        1190:  q   <=  32'b10111111110100010000111110101011 ;
        1191:  q   <=  32'b00111110110101001011100001011000 ;
        1192:  q   <=  32'b10111111001001111001111011101110 ;
        1193:  q   <=  32'b10111110100101111011101011110111 ;
        1194:  q   <=  32'b10111111101111111001101100001001 ;
        1195:  q   <=  32'b10111111011001111010001100111010 ;
        1196:  q   <=  32'b10111110110011101111000011100010 ;
        1197:  q   <=  32'b10111111001110011100110111101000 ;
        1198:  q   <=  32'b10111111010111011101000111110110 ;
        1199:  q   <=  32'b10111110110101111111110001001101 ;
        1200:  q   <=  32'b10111111011100010101001010010100 ;
        1201:  q   <=  32'b00111111101010111100001011011000 ;
        1202:  q   <=  32'b10111111011111010000101000001110 ;
        1203:  q   <=  32'b00111111111010001011001001011000 ;
        1204:  q   <=  32'b10111110101111111011011000100111 ;
        1205:  q   <=  32'b10111111101110011101001010100011 ;
        1206:  q   <=  32'b10111111000111100110000111101110 ;
        1207:  q   <=  32'b00111111011011110011101101110100 ;
        1208:  q   <=  32'b00111111100001110010100010110000 ;
        1209:  q   <=  32'b00111110001001000001001010011110 ;
        1210:  q   <=  32'b00111110100100110010011000100010 ;
        1211:  q   <=  32'b00111111001000100000011000011001 ;
        1212:  q   <=  32'b10111111101110101100000111100010 ;
        1213:  q   <=  32'b10111111000101001110101011101101 ;
        1214:  q   <=  32'b10111111111010100100001001010101 ;
        1215:  q   <=  32'b10111110111001011111000011010110 ;
        1216:  q   <=  32'b00111111011100110000001110101010 ;
        1217:  q   <=  32'b00111111001101111010101000111101 ;
        1218:  q   <=  32'b01000000000100100110101111001000 ;
        1219:  q   <=  32'b00111110001010101011101010101000 ;
        1220:  q   <=  32'b11000000000010100000001111110001 ;
        1221:  q   <=  32'b00111111110110000011111000111100 ;
        1222:  q   <=  32'b00111111101001000010000111000110 ;
        1223:  q   <=  32'b10111111000101010010011101001101 ;
        1224:  q   <=  32'b00111110011000111111010100001100 ;
        1225:  q   <=  32'b00111111010001111000101000100001 ;
        1226:  q   <=  32'b00111110110001001111100001010110 ;
        1227:  q   <=  32'b00111111001100100100010100011010 ;
        1228:  q   <=  32'b10111101111001101101011101101010 ;
        1229:  q   <=  32'b10111101000111110000010110011001 ;
        1230:  q   <=  32'b00111101101101000110011111001111 ;
        1231:  q   <=  32'b10111111010010100010011011100100 ;
        1232:  q   <=  32'b00111111101101100010001110010010 ;
        1233:  q   <=  32'b00111011110011110111101000000100 ;
        1234:  q   <=  32'b00111111001011111011110100110101 ;
        1235:  q   <=  32'b10111111010110101101110011101110 ;
        1236:  q   <=  32'b10111111100010011010000101001111 ;
        1237:  q   <=  32'b10111101101110100100110100001001 ;
        1238:  q   <=  32'b10111110100000010110101101001111 ;
        1239:  q   <=  32'b00111111100110001110111111111100 ;
        1240:  q   <=  32'b00111111000110110010011011111101 ;
        1241:  q   <=  32'b00111111000010100101111100100111 ;
        1242:  q   <=  32'b10111111101110001111001111000110 ;
        1243:  q   <=  32'b10111111011101111011101011001000 ;
        1244:  q   <=  32'b00111110010011101110011010001011 ;
        1245:  q   <=  32'b10111110101100100001110100001111 ;
        1246:  q   <=  32'b00111111101001010010000110011010 ;
        1247:  q   <=  32'b00111111101010111010101011101101 ;
        1248:  q   <=  32'b10111111000101001010111100101000 ;
        1249:  q   <=  32'b00111111011000000000100011100011 ;
        1250:  q   <=  32'b00111111101100101001111000011010 ;
        1251:  q   <=  32'b00111110101001000101100000101100 ;
        1252:  q   <=  32'b00111111110011111100101011111111 ;
        1253:  q   <=  32'b00111111100001111111110111010000 ;
        1254:  q   <=  32'b00111110010110110011111001100111 ;
        1255:  q   <=  32'b00111111011000000111011000101100 ;
        1256:  q   <=  32'b00111110010001110001001010100001 ;
        1257:  q   <=  32'b10111110110101000110110010111110 ;
        1258:  q   <=  32'b00111110101101111000011111100111 ;
        1259:  q   <=  32'b00111101000101000101111000111000 ;
        1260:  q   <=  32'b10111110101110101011000011101111 ;
        1261:  q   <=  32'b00111111111000101011000011000100 ;
        1262:  q   <=  32'b00111110011000101001010101101000 ;
        1263:  q   <=  32'b01000000001011101011111010000001 ;
        1264:  q   <=  32'b10111110100101111010001011111101 ;
        1265:  q   <=  32'b00111111000100000111010110101100 ;
        1266:  q   <=  32'b00111111110010101001001101010000 ;
        1267:  q   <=  32'b01000000001011101010101110110100 ;
        1268:  q   <=  32'b00111110100110110110110011000111 ;
        1269:  q   <=  32'b10111111010010100100111001100001 ;
        1270:  q   <=  32'b00111111010011011010101001010011 ;
        1271:  q   <=  32'b10111111101010001111001010010010 ;
        1272:  q   <=  32'b10111110100011000011010110000010 ;
        1273:  q   <=  32'b00111110100010110011001000100100 ;
        1274:  q   <=  32'b00111111101111101010100110110000 ;
        1275:  q   <=  32'b00111111101101111111010001000000 ;
        1276:  q   <=  32'b10111100111000011100100001110000 ;
        1277:  q   <=  32'b00111111011011001000011011000011 ;
        1278:  q   <=  32'b10111110101001000111111011011110 ;
        1279:  q   <=  32'b00111111001010010011111101111011 ;
        1280:  q   <=  32'b00111111111101010010100001011010 ;
        1281:  q   <=  32'b00111110001000001000010110010111 ;
        1282:  q   <=  32'b10111110100110011101111111101010 ;
        1283:  q   <=  32'b10111111000000000000001001000111 ;
        1284:  q   <=  32'b00111111001101110110101010101011 ;
        1285:  q   <=  32'b00111111101010110010110001000110 ;
        1286:  q   <=  32'b01000000000010000000101100100011 ;
        1287:  q   <=  32'b00111101010111010101111100011100 ;
        1288:  q   <=  32'b00111110001001101111001011100011 ;
        1289:  q   <=  32'b10111111001000011111100100010001 ;
        1290:  q   <=  32'b00111111110011100101010110111100 ;
        1291:  q   <=  32'b10111101100110101000010011011100 ;
        1292:  q   <=  32'b10111110111100100100110000100011 ;
        1293:  q   <=  32'b01000000000010111100101010011001 ;
        1294:  q   <=  32'b00111111010011110101010001011110 ;
        1295:  q   <=  32'b00111111001101110110001000111101 ;
        1296:  q   <=  32'b10111111100000001011011010001110 ;
        1297:  q   <=  32'b00111110110111100011001101111110 ;
        1298:  q   <=  32'b00111111000001010010100000100001 ;
        1299:  q   <=  32'b10111111100010111100111010101011 ;
        1300:  q   <=  32'b10111110011001110011011010101001 ;
        1301:  q   <=  32'b10111110110011110101000111101000 ;
        1302:  q   <=  32'b00111111000001110010000111001000 ;
        1303:  q   <=  32'b10111111100000001110010000101000 ;
        1304:  q   <=  32'b00111111100010110110010100111010 ;
        1305:  q   <=  32'b00111111111001000111011011000110 ;
        1306:  q   <=  32'b10111110100110111000010110110110 ;
        1307:  q   <=  32'b10111100000011100111110001010000 ;
        1308:  q   <=  32'b00111111000000011011001011010101 ;
        1309:  q   <=  32'b00111111100110100000010000101001 ;
        1310:  q   <=  32'b00111111000001011010001011110100 ;
        1311:  q   <=  32'b00111110110010110100100110100000 ;
        1312:  q   <=  32'b10111110111101110011001011111011 ;
        1313:  q   <=  32'b10111110011011010000110110011001 ;
        1314:  q   <=  32'b00111111000111010000011011010000 ;
        1315:  q   <=  32'b00111111110101110110011110100101 ;
        1316:  q   <=  32'b00111111000100011000001000111101 ;
        1317:  q   <=  32'b10111111100110100101111100101010 ;
        1318:  q   <=  32'b00111110110111011011101000010111 ;
        1319:  q   <=  32'b10111101101111001010100111001101 ;
        1320:  q   <=  32'b10111110011110011110100110001001 ;
        1321:  q   <=  32'b10111110011000000111001011111110 ;
        1322:  q   <=  32'b10111111011000010011100001100100 ;
        1323:  q   <=  32'b10111110101001000100000001110110 ;
        1324:  q   <=  32'b10111111010010001100111101110000 ;
        1325:  q   <=  32'b10111110101110101101110001011110 ;
        1326:  q   <=  32'b00111101111100000010101110001101 ;
        1327:  q   <=  32'b00111110001100101000011000011010 ;
        1328:  q   <=  32'b10111110010111001101010100001000 ;
        1329:  q   <=  32'b10111110000111000100011000101111 ;
        1330:  q   <=  32'b00111101000010011111110010101000 ;
        1331:  q   <=  32'b00111110111010101010001111110111 ;
        1332:  q   <=  32'b00111111101001000000110001111101 ;
        1333:  q   <=  32'b00111111000111101011111000111000 ;
        1334:  q   <=  32'b10111110100100101100011011101010 ;
        1335:  q   <=  32'b00111111000110010001011110001110 ;
        1336:  q   <=  32'b10111110011110110110110011101010 ;
        1337:  q   <=  32'b10111111111000111110111100110010 ;
        1338:  q   <=  32'b11000000000101100011100100101010 ;
        1339:  q   <=  32'b10111111110110110101011100010111 ;
        1340:  q   <=  32'b10111110011100101101000101111101 ;
        1341:  q   <=  32'b10111111000111101001111111001100 ;
        1342:  q   <=  32'b10111111001110000101110001101110 ;
        1343:  q   <=  32'b00111101001001101000100000100010 ;
        1344:  q   <=  32'b10111111001010001011001100000001 ;
        1345:  q   <=  32'b10111111001000010110100101101110 ;
        1346:  q   <=  32'b00111111000111000001000001100011 ;
        1347:  q   <=  32'b00111111010010000100011100011010 ;
        1348:  q   <=  32'b01000000000110111111000011111111 ;
        1349:  q   <=  32'b00111110100110101101010100100101 ;
        1350:  q   <=  32'b00111101011011101110000011001100 ;
        1351:  q   <=  32'b10111111000100101111101001110001 ;
        1352:  q   <=  32'b10111110010001111110010111000010 ;
        1353:  q   <=  32'b10111101010011101111100111100010 ;
        1354:  q   <=  32'b10111111111000001011110100111100 ;
        1355:  q   <=  32'b10111110100000111100010001100000 ;
        1356:  q   <=  32'b00111111001111111110000111111010 ;
        1357:  q   <=  32'b10111111000100100001110110011100 ;
        1358:  q   <=  32'b00111110111111010000110000101000 ;
        1359:  q   <=  32'b00111111011111011100111100001010 ;
        1360:  q   <=  32'b00111111100010011101111110111010 ;
        1361:  q   <=  32'b00111111010001101101111100011010 ;
        1362:  q   <=  32'b11000000000100001010000100111001 ;
        1363:  q   <=  32'b10111111000100000111101011111101 ;
        1364:  q   <=  32'b00111111011001101100100000100100 ;
        1365:  q   <=  32'b00111110110010100001001011101001 ;
        1366:  q   <=  32'b00111011100111110001000111011011 ;
        1367:  q   <=  32'b00111110110111111011001111001100 ;
        1368:  q   <=  32'b00111111100100001010011000111001 ;
        1369:  q   <=  32'b00111110000111010111011000010011 ;
        1370:  q   <=  32'b10111111010000100011010101100011 ;
        1371:  q   <=  32'b10111110001110000111110010101100 ;
        1372:  q   <=  32'b10111110010101001100011011001011 ;
        1373:  q   <=  32'b00111111011001011001000100011001 ;
        1374:  q   <=  32'b00111110110100110001100111111110 ;
        1375:  q   <=  32'b00111111000011000010101001000000 ;
        1376:  q   <=  32'b00111110000101110110001000010001 ;
        1377:  q   <=  32'b10111110101110010111101100010100 ;
        1378:  q   <=  32'b00111101011110100110111101001011 ;
        1379:  q   <=  32'b00111110010111011110100000001111 ;
        1380:  q   <=  32'b10111111101100101111010110101100 ;
        1381:  q   <=  32'b00111110001101110010100111001011 ;
        1382:  q   <=  32'b00111111011011010111011000101000 ;
        1383:  q   <=  32'b10111101111000011010010011111000 ;
        1384:  q   <=  32'b00111111110010010100010001010101 ;
        1385:  q   <=  32'b00111111000011110111110001010000 ;
        1386:  q   <=  32'b10111110110101110011011101101000 ;
        1387:  q   <=  32'b10111110000111011010001111011100 ;
        1388:  q   <=  32'b10111110100011001110011011010100 ;
        1389:  q   <=  32'b00111110011101101110100001000111 ;
        1390:  q   <=  32'b00111111010000010011001100100000 ;
        1391:  q   <=  32'b10111110100101010111010100110110 ;
        1392:  q   <=  32'b00111110111010101011100101011010 ;
        1393:  q   <=  32'b00111111111000001010110101001100 ;
        1394:  q   <=  32'b00111111011011100111011000101010 ;
        1395:  q   <=  32'b00111111010100110100010010000111 ;
        1396:  q   <=  32'b10111111010100001001011100110011 ;
        1397:  q   <=  32'b10111111000010001100000110011010 ;
        1398:  q   <=  32'b00111110011110000101111101110110 ;
        1399:  q   <=  32'b10111101110011100010000010000011 ;
        1400:  q   <=  32'b10111111110100000000000110010110 ;
        1401:  q   <=  32'b10111111110000011101100010011110 ;
        1402:  q   <=  32'b00111111100000110101101000101100 ;
        1403:  q   <=  32'b10111111010000100001010010100100 ;
        1404:  q   <=  32'b01000000000001010000001110011001 ;
        1405:  q   <=  32'b11000000000011100011010100000111 ;
        1406:  q   <=  32'b00111110111001011100010001011000 ;
        1407:  q   <=  32'b00111010001001000010000111100100 ;
        1408:  q   <=  32'b10111111010000011001100011100110 ;
        1409:  q   <=  32'b00111110110011110000001110101001 ;
        1410:  q   <=  32'b10111111010010110011100111110001 ;
        1411:  q   <=  32'b00111111010111000001101011000000 ;
        1412:  q   <=  32'b00111101100010001111001010111001 ;
        1413:  q   <=  32'b10111111110100011101011101110010 ;
        1414:  q   <=  32'b11000000000110110010111100011010 ;
        1415:  q   <=  32'b10111110100100010101001000100111 ;
        1416:  q   <=  32'b00111111100100101010100111000111 ;
        1417:  q   <=  32'b00111110001110011000010001110001 ;
        1418:  q   <=  32'b00111101010111100011010101111100 ;
        1419:  q   <=  32'b00111111001100000001000010011111 ;
        1420:  q   <=  32'b10111111101100100101101100101011 ;
        1421:  q   <=  32'b00111111101101100111001001100010 ;
        1422:  q   <=  32'b10111111011001001101001101101101 ;
        1423:  q   <=  32'b00111101000110101010111100101000 ;
        1424:  q   <=  32'b10111110101110100010010111000000 ;
        1425:  q   <=  32'b00111110000110010010010101010101 ;
        1426:  q   <=  32'b10111111111110001110010111111000 ;
        1427:  q   <=  32'b00111111110000110000111011111100 ;
        1428:  q   <=  32'b00111111000010111011101000110111 ;
        1429:  q   <=  32'b01000000000000001010001010100110 ;
        1430:  q   <=  32'b00111111101101010101010101110110 ;
        1431:  q   <=  32'b00111100001111000001100101100110 ;
        1432:  q   <=  32'b10111111011100000110010110001001 ;
        1433:  q   <=  32'b10111111110111101001010010001100 ;
        1434:  q   <=  32'b00111100100010110000011010110100 ;
        1435:  q   <=  32'b00111110011000000110101100111101 ;
        1436:  q   <=  32'b00111111100001011101110101110011 ;
        1437:  q   <=  32'b10111111011100110111001110011001 ;
        1438:  q   <=  32'b00111111010010110111011111011000 ;
        1439:  q   <=  32'b00111101100100100100100111001010 ;
        1440:  q   <=  32'b10111111010001100001000001011000 ;
        1441:  q   <=  32'b00111111010001100010111101111000 ;
        1442:  q   <=  32'b00111110100010000000001111100101 ;
        1443:  q   <=  32'b10111110011100001011111110000001 ;
        1444:  q   <=  32'b00111111111100000100101100011100 ;
        1445:  q   <=  32'b00111111000110111111011100011101 ;
        1446:  q   <=  32'b10111101111000011101011101000101 ;
        1447:  q   <=  32'b00111110100011100000111011100111 ;
        1448:  q   <=  32'b00111101101100100100010100100000 ;
        1449:  q   <=  32'b00111110001100011100001001100000 ;
        1450:  q   <=  32'b00111110111010000011110100011001 ;
        1451:  q   <=  32'b10111111000110101000000000101000 ;
        1452:  q   <=  32'b10111111010011000000100111000010 ;
        1453:  q   <=  32'b00111110101110001010011011111000 ;
        1454:  q   <=  32'b00111111111100010100101010101111 ;
        1455:  q   <=  32'b10111110100111010001011111000000 ;
        1456:  q   <=  32'b10111111100000011010000011110000 ;
        1457:  q   <=  32'b10111110011101000100010101000110 ;
        1458:  q   <=  32'b10111110111101111101000011001010 ;
        1459:  q   <=  32'b10111110101001111001100110110011 ;
        1460:  q   <=  32'b00111110111100110111011100010111 ;
        1461:  q   <=  32'b10111110000001010010000000000000 ;
        1462:  q   <=  32'b10111111000110000010011110001001 ;
        1463:  q   <=  32'b10111110111000110011010101101010 ;
        1464:  q   <=  32'b10111111101010010100100010100110 ;
        1465:  q   <=  32'b10111111010111000000100110010100 ;
        1466:  q   <=  32'b10111111101101001101110100111000 ;
        1467:  q   <=  32'b10111111000001000001011110100110 ;
        1468:  q   <=  32'b10111111100010101110010001111110 ;
        1469:  q   <=  32'b10111111001101010000100001011000 ;
        1470:  q   <=  32'b10111110100110100111001001110110 ;
        1471:  q   <=  32'b10111111100110011010100000001000 ;
        1472:  q   <=  32'b10111100100111101001110110011101 ;
        1473:  q   <=  32'b00111110101011100100010100001100 ;
        1474:  q   <=  32'b10111111011101101001011001001110 ;
        1475:  q   <=  32'b00111111100011101001010100000011 ;
        1476:  q   <=  32'b10111111110010110000010110000000 ;
        1477:  q   <=  32'b10111110110010001001100101001111 ;
        1478:  q   <=  32'b10111111101111100000101000110010 ;
        1479:  q   <=  32'b10111110101100000111001011111000 ;
        1480:  q   <=  32'b10111111101010010111011000010011 ;
        1481:  q   <=  32'b10111111000100110010100001100010 ;
        1482:  q   <=  32'b10111111001111011001111011110100 ;
        1483:  q   <=  32'b10111111100101111010111000100100 ;
        1484:  q   <=  32'b11000000000001000010011010101010 ;
        1485:  q   <=  32'b00111111000100001010011111000010 ;
        1486:  q   <=  32'b01000000000000000000001001010101 ;
        1487:  q   <=  32'b01000000000011100100101100000000 ;
        1488:  q   <=  32'b10111110111110111111111010110011 ;
        1489:  q   <=  32'b10111101001111000110110110010010 ;
        1490:  q   <=  32'b10111110111011100111011001100100 ;
        1491:  q   <=  32'b00111101100110111000101001010011 ;
        1492:  q   <=  32'b10111111011010110011010001111100 ;
        1493:  q   <=  32'b10111111111101011011000100010100 ;
        1494:  q   <=  32'b10111101000101010100010101100111 ;
        1495:  q   <=  32'b10111111100111001101000011101011 ;
        1496:  q   <=  32'b10111111111100111000001011110111 ;
        1497:  q   <=  32'b01000000000101111111001110110000 ;
        1498:  q   <=  32'b10111110011011101111001000101101 ;
        1499:  q   <=  32'b00111110110011101100100101110100 ;
        1500:  q   <=  32'b00111111100110001010001011001111 ;
        1501:  q   <=  32'b10111111110101111010011000101101 ;
        1502:  q   <=  32'b00111110110100111000100000110100 ;
        1503:  q   <=  32'b00111111000000000111001001011111 ;
        1504:  q   <=  32'b00111101101010100001110110100011 ;
        1505:  q   <=  32'b00111110001000011001010111010000 ;
        1506:  q   <=  32'b10111111000001110010011100111101 ;
        1507:  q   <=  32'b00111111001110010001101010000001 ;
        1508:  q   <=  32'b10111111010110011001010111000110 ;
        1509:  q   <=  32'b10111111010010111101111111010011 ;
        1510:  q   <=  32'b00111111001110011010111110111001 ;
        1511:  q   <=  32'b00111111110101111110000010110000 ;
        1512:  q   <=  32'b10111110110001011101010101110100 ;
        1513:  q   <=  32'b10111111000000010100110011010001 ;
        1514:  q   <=  32'b00111110110100001110111100001111 ;
        1515:  q   <=  32'b00111111100010010100001011110111 ;
        1516:  q   <=  32'b00111111011101111100110110111010 ;
        1517:  q   <=  32'b00111110100010100101000010000011 ;
        1518:  q   <=  32'b10111111001000100110100001110111 ;
        1519:  q   <=  32'b00111111001000010011100000101000 ;
        1520:  q   <=  32'b10111101101000100100010101001110 ;
        1521:  q   <=  32'b00111111101100000011111111011110 ;
        1522:  q   <=  32'b10111111101101000100000001001110 ;
        1523:  q   <=  32'b00111110000100001001111100001001 ;
        1524:  q   <=  32'b00111111101001010001010110000110 ;
        1525:  q   <=  32'b10111110111111010110100001001010 ;
        1526:  q   <=  32'b10111111000111111111010010000111 ;
        1527:  q   <=  32'b10111111011011110000001010101000 ;
        1528:  q   <=  32'b10111110100011101011010100001000 ;
        1529:  q   <=  32'b10111110010011010101011001101010 ;
        1530:  q   <=  32'b00111110000011000000010111100000 ;
        1531:  q   <=  32'b10111111011000100010001100100110 ;
        1532:  q   <=  32'b00111101101010010000100110100100 ;
        1533:  q   <=  32'b10111111000110101001011110001011 ;
        1534:  q   <=  32'b10111110101111001100100111110011 ;
        1535:  q   <=  32'b10111111010101101001001001010110 ;
        1536:  q   <=  32'b10111110100100001010000010010001 ;
        1537:  q   <=  32'b01000000011001000111100010110110 ;
        1538:  q   <=  32'b01000000010110100001010100000010 ;
        1539:  q   <=  32'b00111111100100101100111000110100 ;
        1540:  q   <=  32'b00111111010010011000100110110101 ;
        1541:  q   <=  32'b10111111101000111001101000000001 ;
        1542:  q   <=  32'b10111111000101011010011111100100 ;
        1543:  q   <=  32'b10111111000111101001000101011110 ;
        1544:  q   <=  32'b00111111000010010000100101111101 ;
        1545:  q   <=  32'b00111110111101110100101000010100 ;
        1546:  q   <=  32'b00111101110111100010100000101111 ;
        1547:  q   <=  32'b10111110101011100011100111001100 ;
        1548:  q   <=  32'b10111111011011010000010001100110 ;
        1549:  q   <=  32'b00111011101011100110000110010001 ;
        1550:  q   <=  32'b00111111100100011100111110100110 ;
        1551:  q   <=  32'b00111110110110101100111100010111 ;
        1552:  q   <=  32'b00111110001110010110000001111101 ;
        1553:  q   <=  32'b00111111001010000101000010010111 ;
        1554:  q   <=  32'b00111111000101011001000100011110 ;
        1555:  q   <=  32'b10111111110011101110011111100000 ;
        1556:  q   <=  32'b00111100100110011100110010101011 ;
        1557:  q   <=  32'b10111110110110100001011110000111 ;
        1558:  q   <=  32'b11000000000000100010110110000000 ;
        1559:  q   <=  32'b10111111101010100000111000000010 ;
        1560:  q   <=  32'b10111110101000111100100000001100 ;
        1561:  q   <=  32'b00111111010100110100111101101001 ;
        1562:  q   <=  32'b10111110011010101100101110111011 ;
        1563:  q   <=  32'b00111110100001100100010110111101 ;
        1564:  q   <=  32'b10111111011001011110000111111100 ;
        1565:  q   <=  32'b11000000000010100001000100111111 ;
        1566:  q   <=  32'b00111101110000000101011101101101 ;
        1567:  q   <=  32'b10111111011100111000000010100000 ;
        1568:  q   <=  32'b00111111100101100001011101101101 ;
        1569:  q   <=  32'b00111111110111100001011110011111 ;
        1570:  q   <=  32'b10111110101111100100111011110001 ;
        1571:  q   <=  32'b00111111100110001010111111000101 ;
        1572:  q   <=  32'b00111111011101000010001001000110 ;
        1573:  q   <=  32'b10111111101101010010000000101101 ;
        1574:  q   <=  32'b10111101000010001010000010100010 ;
        1575:  q   <=  32'b00111110100001011011000100111010 ;
        1576:  q   <=  32'b00111111000001011110001011111000 ;
        1577:  q   <=  32'b00111111001011010100000111100111 ;
        1578:  q   <=  32'b00111111001011001010010100110001 ;
        1579:  q   <=  32'b00111111001011011010101110001101 ;
        1580:  q   <=  32'b10111110101000000000101001110010 ;
        1581:  q   <=  32'b00111110110000100010110000111101 ;
        1582:  q   <=  32'b11000000000100000010111101111100 ;
        1583:  q   <=  32'b10111111100101011000110010000100 ;
        1584:  q   <=  32'b00111111100110011101101000000010 ;
        1585:  q   <=  32'b10111111001010010010011000101010 ;
        1586:  q   <=  32'b00111110101001111011010111010001 ;
        1587:  q   <=  32'b00111111110000010000101001001110 ;
        1588:  q   <=  32'b10111111011000111000111110001001 ;
        1589:  q   <=  32'b10111111011101011001001110101101 ;
        1590:  q   <=  32'b10111110111111000100010110110100 ;
        1591:  q   <=  32'b00111110111000011101001000101010 ;
        1592:  q   <=  32'b10111110010100011010110110111000 ;
        1593:  q   <=  32'b10111111011110100101000110001110 ;
        1594:  q   <=  32'b10111111110010010101011001010000 ;
        1595:  q   <=  32'b10111110101111011001001011101100 ;
        1596:  q   <=  32'b10111110011000100111001111110101 ;
        1597:  q   <=  32'b10111111000010010000001110110101 ;
        1598:  q   <=  32'b10111110100001100010000100110111 ;
        1599:  q   <=  32'b10111111100011000011011010001110 ;
        1600:  q   <=  32'b00111111000011001001101010010000 ;
        1601:  q   <=  32'b11000000000010110010110011111011 ;
        1602:  q   <=  32'b00111110000101000001010111011100 ;
        1603:  q   <=  32'b00111111001010110100010111000110 ;
        1604:  q   <=  32'b10111111010110010100110011011110 ;
        1605:  q   <=  32'b10111101011010011101011101010100 ;
        1606:  q   <=  32'b00111110100101010110010100000010 ;
        1607:  q   <=  32'b10111111000111010101011110100100 ;
        1608:  q   <=  32'b10111100010111111000011110101110 ;
        1609:  q   <=  32'b00111110110100110000000010001010 ;
        1610:  q   <=  32'b10111111011011111110100100001001 ;
        1611:  q   <=  32'b00111111010101011100110011011001 ;
        1612:  q   <=  32'b00111111100011000001100111010110 ;
        1613:  q   <=  32'b00111110101001000111000111001101 ;
        1614:  q   <=  32'b00111100011101111001101111010110 ;
        1615:  q   <=  32'b10111111100101010000111000010111 ;
        1616:  q   <=  32'b00111110111111010101101111000100 ;
        1617:  q   <=  32'b10111111100110111010000011110000 ;
        1618:  q   <=  32'b00111111110010111001111011110000 ;
        1619:  q   <=  32'b00111111000001101100011100010001 ;
        1620:  q   <=  32'b00111110100001111001011001001101 ;
        1621:  q   <=  32'b10111110110010011000010110101001 ;
        1622:  q   <=  32'b11000000000010110100100010101001 ;
        1623:  q   <=  32'b10111111100110010000101100110100 ;
        1624:  q   <=  32'b00111110101110110000110001010010 ;
        1625:  q   <=  32'b01000000000110100110010101110111 ;
        1626:  q   <=  32'b00111111001111011000000011010111 ;
        1627:  q   <=  32'b00111110100111101001011100010100 ;
        1628:  q   <=  32'b10111111000010101011111110101100 ;
        1629:  q   <=  32'b00111101111110100110111110011011 ;
        1630:  q   <=  32'b00111111011101100101011111110000 ;
        1631:  q   <=  32'b10111110100000100000100011111101 ;
        1632:  q   <=  32'b00111111111100100010010100001111 ;
        1633:  q   <=  32'b10111111100111000011000101001001 ;
        1634:  q   <=  32'b10111110110000001010001000100111 ;
        1635:  q   <=  32'b00111101010101101011111111110010 ;
        1636:  q   <=  32'b10111111111110100001101001111111 ;
        1637:  q   <=  32'b00111111000100001011111101100111 ;
        1638:  q   <=  32'b00111101100111110101001010110011 ;
        1639:  q   <=  32'b00111101101001010100011010101010 ;
        1640:  q   <=  32'b00111111010010110111000111111000 ;
        1641:  q   <=  32'b00111111100001011001011110011001 ;
        1642:  q   <=  32'b00111111010011010101101111111001 ;
        1643:  q   <=  32'b10111110111100000000100110111111 ;
        1644:  q   <=  32'b10111101001111101101011110100101 ;
        1645:  q   <=  32'b00111110101101001111011111001011 ;
        1646:  q   <=  32'b10111111101000001101111011010111 ;
        1647:  q   <=  32'b10111111100001001001110010101101 ;
        1648:  q   <=  32'b10111110110110101001101011011010 ;
        1649:  q   <=  32'b00111101100111110001000011000001 ;
        1650:  q   <=  32'b00111111111001010011110100110011 ;
        1651:  q   <=  32'b00111111010011000001100101101111 ;
        1652:  q   <=  32'b10111110111000101000111101110101 ;
        1653:  q   <=  32'b10111111001000010000110000011101 ;
        1654:  q   <=  32'b00111111110001000101001101101111 ;
        1655:  q   <=  32'b01000000001011101111001001010011 ;
        1656:  q   <=  32'b00111110001010110111010100100110 ;
        1657:  q   <=  32'b10111110111101010010110111010000 ;
        1658:  q   <=  32'b10111111101101001101000111010111 ;
        1659:  q   <=  32'b00111111011110011001100011010001 ;
        1660:  q   <=  32'b00111110100101000101011000001011 ;
        1661:  q   <=  32'b00111111100101010010110000011000 ;
        1662:  q   <=  32'b10111111011010001010000011101110 ;
        1663:  q   <=  32'b00111110011101100101100101001101 ;
        1664:  q   <=  32'b10111111001001110110111110010100 ;
        1665:  q   <=  32'b00111111101000110011000110110101 ;
        1666:  q   <=  32'b10111111000011010001101011010011 ;
        1667:  q   <=  32'b10111101101100110000001101101011 ;
        1668:  q   <=  32'b10111110101100100001010110000001 ;
        1669:  q   <=  32'b00111111011111100111010001010100 ;
        1670:  q   <=  32'b00111110110110110101101111111100 ;
        1671:  q   <=  32'b10111111100000001000100100100100 ;
        1672:  q   <=  32'b10111111001000011111011111010101 ;
        1673:  q   <=  32'b10111111100001011101100111010011 ;
        1674:  q   <=  32'b00111111000000010111011000000011 ;
        1675:  q   <=  32'b00111110101010011111010111010110 ;
        1676:  q   <=  32'b10111111110100010101010100110010 ;
        1677:  q   <=  32'b10111111111101000001001101010111 ;
        1678:  q   <=  32'b10111101001001010111100100100001 ;
        1679:  q   <=  32'b00111111001100100111101101000011 ;
        1680:  q   <=  32'b00111110001011001101101010010101 ;
        1681:  q   <=  32'b10111111110001011001101100011110 ;
        1682:  q   <=  32'b10111111110001101010000101110101 ;
        1683:  q   <=  32'b00111111010111011111100011001111 ;
        1684:  q   <=  32'b10111110000101001101110010101000 ;
        1685:  q   <=  32'b10111110110001011100000101110111 ;
        1686:  q   <=  32'b00111111101010000111100101100000 ;
        1687:  q   <=  32'b10111111010010111110010100010100 ;
        1688:  q   <=  32'b00111110000010101011000100100100 ;
        1689:  q   <=  32'b00111110110101011110101010111001 ;
        1690:  q   <=  32'b00111111010100011110001110100001 ;
        1691:  q   <=  32'b10111111010110101011011011100111 ;
        1692:  q   <=  32'b00111110101101101111001001110110 ;
        1693:  q   <=  32'b01000000001011111110011011100000 ;
        1694:  q   <=  32'b10111111110000011010100100111010 ;
        1695:  q   <=  32'b00111110110111100011001001111111 ;
        1696:  q   <=  32'b10111110011010110100100000111011 ;
        1697:  q   <=  32'b10111111010100111011101111101110 ;
        1698:  q   <=  32'b10111111010101001111110011010000 ;
        1699:  q   <=  32'b00111110111111101110110010101110 ;
        1700:  q   <=  32'b01000000000101000011001100110111 ;
        1701:  q   <=  32'b10111111010010110011100000101001 ;
        1702:  q   <=  32'b00111111000010100111110001010011 ;
        1703:  q   <=  32'b10111111000011110001111010100101 ;
        1704:  q   <=  32'b00111111111111010000000000011101 ;
        1705:  q   <=  32'b00111111000010110110111011011100 ;
        1706:  q   <=  32'b10111110000011010011011100011101 ;
        1707:  q   <=  32'b00111111000111101011000000101011 ;
        1708:  q   <=  32'b10111011101101101110111111001000 ;
        1709:  q   <=  32'b00111111100011011011100010110100 ;
        1710:  q   <=  32'b10111110001111100000101101010101 ;
        1711:  q   <=  32'b10111111100011111000101010011110 ;
        1712:  q   <=  32'b00111110011111000101110101000011 ;
        1713:  q   <=  32'b00111111110001111101000000010001 ;
        1714:  q   <=  32'b10111111100110010010101011100110 ;
        1715:  q   <=  32'b10111110011110000010100101011100 ;
        1716:  q   <=  32'b00111111100000001001111000110101 ;
        1717:  q   <=  32'b10111111111101011100011010101110 ;
        1718:  q   <=  32'b00111111001000000001110100110110 ;
        1719:  q   <=  32'b00111111010000001100001000000011 ;
        1720:  q   <=  32'b00111110010110101001101101110111 ;
        1721:  q   <=  32'b10111111010001010010111000001111 ;
        1722:  q   <=  32'b10111011111010011100100111001101 ;
        1723:  q   <=  32'b00111101101111101101100010010011 ;
        1724:  q   <=  32'b00111111011011110110110010011111 ;
        1725:  q   <=  32'b00111111001010011101110001001111 ;
        1726:  q   <=  32'b10111110101100110101000110110010 ;
        1727:  q   <=  32'b00111111110011110101100000100100 ;
        1728:  q   <=  32'b10111101010100000011011001011101 ;
        1729:  q   <=  32'b10111111010100000000110011101010 ;
        1730:  q   <=  32'b10111110111000000111100010010011 ;
        1731:  q   <=  32'b00111111010110111100110111011101 ;
        1732:  q   <=  32'b00111110010001111110011010101111 ;
        1733:  q   <=  32'b00111111011000111000110001111000 ;
        1734:  q   <=  32'b00111101100011011100010000101011 ;
        1735:  q   <=  32'b01000000000111110010100000010100 ;
        1736:  q   <=  32'b10111111110101010011001111001011 ;
        1737:  q   <=  32'b10111110110101001111010010000001 ;
        1738:  q   <=  32'b10111101101011000111110111110011 ;
        1739:  q   <=  32'b00111101101101101100100110111001 ;
        1740:  q   <=  32'b00111111101110100110001100001000 ;
        1741:  q   <=  32'b00111110011000001011100001101100 ;
        1742:  q   <=  32'b10111101111010110100010011000011 ;
        1743:  q   <=  32'b00111101100011000111111101110011 ;
        1744:  q   <=  32'b00111111010000000110000111110111 ;
        1745:  q   <=  32'b10111111001100000111111001001010 ;
        1746:  q   <=  32'b00111110111001101101000100001001 ;
        1747:  q   <=  32'b10111111110010000101001010111010 ;
        1748:  q   <=  32'b10111101101000010101111111000001 ;
        1749:  q   <=  32'b10111111011100010001100101000111 ;
        1750:  q   <=  32'b10111111001001110010000111101110 ;
        1751:  q   <=  32'b00111110100100001010011110101100 ;
        1752:  q   <=  32'b10111111100100000000001010010111 ;
        1753:  q   <=  32'b10111111011111010010110101100111 ;
        1754:  q   <=  32'b10111111110000100000011110101000 ;
        1755:  q   <=  32'b11000000000011101001111111101010 ;
        1756:  q   <=  32'b10111110000110110010100001111111 ;
        1757:  q   <=  32'b00111111100101001101010011001110 ;
        1758:  q   <=  32'b10111110001110100100110110000001 ;
        1759:  q   <=  32'b10111110011011111001000110000100 ;
        1760:  q   <=  32'b10111111100001011111101101100001 ;
        1761:  q   <=  32'b00111111110010101010101000110001 ;
        1762:  q   <=  32'b10111110011111110110011000111011 ;
        1763:  q   <=  32'b00111111101001011010001001101010 ;
        1764:  q   <=  32'b00111110101110010101010101110101 ;
        1765:  q   <=  32'b10111110100001101010111011010001 ;
        1766:  q   <=  32'b00111111100010101000001110110101 ;
        1767:  q   <=  32'b00111111011110111000000011001100 ;
        1768:  q   <=  32'b10111101111001000011110010111011 ;
        1769:  q   <=  32'b00111111101001011110000110110111 ;
        1770:  q   <=  32'b00111111111001000000000101111001 ;
        1771:  q   <=  32'b10111101100001100110000100010111 ;
        1772:  q   <=  32'b10111110100000101110100010011010 ;
        1773:  q   <=  32'b00111110110011110010110010111011 ;
        1774:  q   <=  32'b00111110101101000001100101110110 ;
        1775:  q   <=  32'b00111111010011101011100100001011 ;
        1776:  q   <=  32'b10111110100000101101110011000001 ;
        1777:  q   <=  32'b00111111001101110001000110101001 ;
        1778:  q   <=  32'b00111111100001100011100001101111 ;
        1779:  q   <=  32'b00111110001101011100111101001001 ;
        1780:  q   <=  32'b00111110000111001111101000010001 ;
        1781:  q   <=  32'b10111111101000001000110110110100 ;
        1782:  q   <=  32'b10111111100101100001111001010110 ;
        1783:  q   <=  32'b10111111101110110001000010000110 ;
        1784:  q   <=  32'b10111111100111110100010011010100 ;
        1785:  q   <=  32'b10111110000111101101001001011110 ;
        1786:  q   <=  32'b10111111110011101011010101111110 ;
        1787:  q   <=  32'b01000000000011111011111110001000 ;
        1788:  q   <=  32'b00111111001111010100000110000111 ;
        1789:  q   <=  32'b11000000000001000101010001001101 ;
        1790:  q   <=  32'b10111111100100111100100001010000 ;
        1791:  q   <=  32'b10111101110110111000011101101010 ;
        1792:  q   <=  32'b10111111110110110011111110011111 ;
        1793:  q   <=  32'b10111110111010110111011101001100 ;
        1794:  q   <=  32'b00111111100010111010010111100100 ;
        1795:  q   <=  32'b10111110001001111101000000111001 ;
        1796:  q   <=  32'b10111101100010011011010101011111 ;
        1797:  q   <=  32'b10111111100000000011010000101110 ;
        1798:  q   <=  32'b10111111000011100011111111010100 ;
        1799:  q   <=  32'b10111111101011001111111111001100 ;
        1800:  q   <=  32'b00111110101110100111100111101000 ;
        1801:  q   <=  32'b10111110111001111000011111000001 ;
        1802:  q   <=  32'b00111111010010001000101010101100 ;
        1803:  q   <=  32'b00111111100111100101110111000101 ;
        1804:  q   <=  32'b00111111100010011110000110100001 ;
        1805:  q   <=  32'b10111101000011101011010110010000 ;
        1806:  q   <=  32'b10111111000000010000010101010000 ;
        1807:  q   <=  32'b10111111100111001010110010100111 ;
        1808:  q   <=  32'b00111101111100101011010011100011 ;
        1809:  q   <=  32'b00111111011101011010000000001110 ;
        1810:  q   <=  32'b10111110101011101000111001101111 ;
        1811:  q   <=  32'b10111110001100010111101001011100 ;
        1812:  q   <=  32'b00111111000111011100010111011110 ;
        1813:  q   <=  32'b00111111010111010010100111010001 ;
        1814:  q   <=  32'b10111111101101010101110101110001 ;
        1815:  q   <=  32'b00111110010011001100000000110100 ;
        1816:  q   <=  32'b00111110010010001000011011010101 ;
        1817:  q   <=  32'b10111110000110101100001001110011 ;
        1818:  q   <=  32'b00111111011001001000110110000000 ;
        1819:  q   <=  32'b10111110101110100111011100100010 ;
        1820:  q   <=  32'b10111111010100111000000100011010 ;
        1821:  q   <=  32'b00111110100011010101000101011010 ;
        1822:  q   <=  32'b00111110111010110110101010001101 ;
        1823:  q   <=  32'b10111110010111101011101000010001 ;
        1824:  q   <=  32'b00111111010010111100111010110110 ;
        1825:  q   <=  32'b10111111110000100100111010010000 ;
        1826:  q   <=  32'b10111111100010011001011011100001 ;
        1827:  q   <=  32'b11000000010001001001111001011101 ;
        1828:  q   <=  32'b00111111000001010111101011110001 ;
        1829:  q   <=  32'b10111111011111011011001110111001 ;
        1830:  q   <=  32'b10111110100000011001100110110010 ;
        1831:  q   <=  32'b00111111100000010010111110011010 ;
        1832:  q   <=  32'b00111101010100001111001000000011 ;
        1833:  q   <=  32'b10111110111000011000000001101000 ;
        1834:  q   <=  32'b10111111010110010011010101001010 ;
        1835:  q   <=  32'b10111110011101100010001111000101 ;
        1836:  q   <=  32'b00111111000110100101100110010101 ;
        1837:  q   <=  32'b10111111110000100001010010011001 ;
        1838:  q   <=  32'b10111101100010111111101001001100 ;
        1839:  q   <=  32'b00111111010010000100101011100110 ;
        1840:  q   <=  32'b10111111101101011101101001011000 ;
        1841:  q   <=  32'b00111111001010110101101110000011 ;
        1842:  q   <=  32'b00111111001011101110100010011000 ;
        1843:  q   <=  32'b10111111011000011101001110101101 ;
        1844:  q   <=  32'b10111111110000001001001110111110 ;
        1845:  q   <=  32'b00111110110111011100010001110010 ;
        1846:  q   <=  32'b00111111010011101110100111011000 ;
        1847:  q   <=  32'b00111111000101000011010101000111 ;
        1848:  q   <=  32'b00111111010000110100101000010100 ;
        1849:  q   <=  32'b10111111100101110100111111110000 ;
        1850:  q   <=  32'b00111111000101010111011100001010 ;
        1851:  q   <=  32'b10111111000101000111101110000011 ;
        1852:  q   <=  32'b10111111000011111011010111000010 ;
        1853:  q   <=  32'b10111111110001110010011110011101 ;
        1854:  q   <=  32'b00111111100011001101001110100001 ;
        1855:  q   <=  32'b00111110001100110100001001111011 ;
        1856:  q   <=  32'b00111111100000000111011001010101 ;
        1857:  q   <=  32'b00111111110000010110100010110111 ;
        1858:  q   <=  32'b10111111100100011001000100001100 ;
        1859:  q   <=  32'b00111111001001001001110011011010 ;
        1860:  q   <=  32'b10111100010100010000111110000000 ;
        1861:  q   <=  32'b00111111011010100000110011101100 ;
        1862:  q   <=  32'b00111111100011011100100011101111 ;
        1863:  q   <=  32'b00111111010100100000101001101010 ;
        1864:  q   <=  32'b10111111010100010100111100000010 ;
        1865:  q   <=  32'b10111110000000011000010101010111 ;
        1866:  q   <=  32'b00111110100001110011110110111101 ;
        1867:  q   <=  32'b01000000010010100010010101010010 ;
        1868:  q   <=  32'b00111111100111010000000111001011 ;
        1869:  q   <=  32'b01000000000101001000010101001010 ;
        1870:  q   <=  32'b00111110110101000011100100010000 ;
        1871:  q   <=  32'b00111110010110001110101001011111 ;
        1872:  q   <=  32'b00111111000111001111100010000001 ;
        1873:  q   <=  32'b10111111000001110001110001100100 ;
        1874:  q   <=  32'b00111111100111101110110011001010 ;
        1875:  q   <=  32'b10111110001000010110100111110000 ;
        1876:  q   <=  32'b10111111101011111101001000101110 ;
        1877:  q   <=  32'b00111111010111101110111100111111 ;
        1878:  q   <=  32'b10111111110010001100010110110011 ;
        1879:  q   <=  32'b10111111111011000001000001111010 ;
        1880:  q   <=  32'b00111110100100111010101001110011 ;
        1881:  q   <=  32'b10111111011100110110111011101001 ;
        1882:  q   <=  32'b10111111011010010010010110111101 ;
        1883:  q   <=  32'b10111110001001011101011000000000 ;
        1884:  q   <=  32'b10111110111110100101000101010101 ;
        1885:  q   <=  32'b10111110011001000010000011110111 ;
        1886:  q   <=  32'b00111110100010110100110001001100 ;
        1887:  q   <=  32'b10111111100101011001001001101011 ;
        1888:  q   <=  32'b10111111100111001011001110110101 ;
        1889:  q   <=  32'b11000000000001100101110111011011 ;
        1890:  q   <=  32'b10111110110001111100110111100001 ;
        1891:  q   <=  32'b00111111001010100000111001011110 ;
        1892:  q   <=  32'b10111111001100111100011110010010 ;
        1893:  q   <=  32'b00111111000000000101011100000000 ;
        1894:  q   <=  32'b00111111000010100101001000000000 ;
        1895:  q   <=  32'b00111111011111011010000111011011 ;
        1896:  q   <=  32'b00111111011111010100011111100010 ;
        1897:  q   <=  32'b10111111001100000101011111100101 ;
        1898:  q   <=  32'b10111111010110110101100110110101 ;
        1899:  q   <=  32'b00111101010001100011010010011100 ;
        1900:  q   <=  32'b10111111001010100011001111010101 ;
        1901:  q   <=  32'b00111111101110011111001101110010 ;
        1902:  q   <=  32'b00111111101100001001111011001001 ;
        1903:  q   <=  32'b00111101110000101101011011100010 ;
        1904:  q   <=  32'b10111110110110101011000001100110 ;
        1905:  q   <=  32'b00111111000000101100010001001100 ;
        1906:  q   <=  32'b10111111001010000000000110001100 ;
        1907:  q   <=  32'b10111110000000000000010001100101 ;
        1908:  q   <=  32'b10111111000001111100110010101010 ;
        1909:  q   <=  32'b00111101110110000011110110101110 ;
        1910:  q   <=  32'b00111111100100000110110111001001 ;
        1911:  q   <=  32'b00111111001111100001001100001010 ;
        1912:  q   <=  32'b00111111100100100110000110010110 ;
        1913:  q   <=  32'b10111111011010100010101010110110 ;
        1914:  q   <=  32'b00111110001110000001110111101101 ;
        1915:  q   <=  32'b10111111011110111011110010101110 ;
        1916:  q   <=  32'b00111110110001010000100001000000 ;
        1917:  q   <=  32'b00111110101001101100000111010111 ;
        1918:  q   <=  32'b00111111101001011110110101111111 ;
        1919:  q   <=  32'b00111111100011001011001110001101 ;
        1920:  q   <=  32'b00111111001001110011100110100000 ;
        1921:  q   <=  32'b10111111000000010100110001111101 ;
        1922:  q   <=  32'b10111110111100111011010101110101 ;
        1923:  q   <=  32'b11000000000000110100110011001000 ;
        1924:  q   <=  32'b10111110111001011000100000101100 ;
        1925:  q   <=  32'b10111111110001101000110110011011 ;
        1926:  q   <=  32'b00111111011011100000100100001111 ;
        1927:  q   <=  32'b00111111011001101110010110001001 ;
        1928:  q   <=  32'b00111110000011011001101100111001 ;
        1929:  q   <=  32'b10111110110000011011111010101001 ;
        1930:  q   <=  32'b00111110000100100111111101101111 ;
        1931:  q   <=  32'b00111111110011010111000111101000 ;
        1932:  q   <=  32'b00111111101011001010111111010101 ;
        1933:  q   <=  32'b10111110111001011001101000110100 ;
        1934:  q   <=  32'b00111110001011000111010000000100 ;
        1935:  q   <=  32'b10111111100011110110110001101111 ;
        1936:  q   <=  32'b00111110110011010010110010011001 ;
        1937:  q   <=  32'b00111111001111010011001100110101 ;
        1938:  q   <=  32'b00111111011001100110100101010100 ;
        1939:  q   <=  32'b10111111110000111111111011110101 ;
        1940:  q   <=  32'b00111111000000010010111011010011 ;
        1941:  q   <=  32'b10111111010111010011110100101011 ;
        1942:  q   <=  32'b10111110110000001100101111001111 ;
        1943:  q   <=  32'b00111111010010011011101100001100 ;
        1944:  q   <=  32'b00111110100110001010111001101000 ;
        1945:  q   <=  32'b10111110001001111010101111110000 ;
        1946:  q   <=  32'b00111111000110110101001011010010 ;
        1947:  q   <=  32'b00111111110100010011011101000000 ;
        1948:  q   <=  32'b10111111000111111001110101001000 ;
        1949:  q   <=  32'b10111111101011001101000000010101 ;
        1950:  q   <=  32'b10111111100101001100010001001111 ;
        1951:  q   <=  32'b10111111011100011011110001001000 ;
        1952:  q   <=  32'b10111111001010111101010001111010 ;
        1953:  q   <=  32'b00111111000100111010000101100000 ;
        1954:  q   <=  32'b11000000000001010111110101000001 ;
        1955:  q   <=  32'b00111110011100011010000010000100 ;
        1956:  q   <=  32'b10111111010001110100011010011111 ;
        1957:  q   <=  32'b00111111100011001011111001110010 ;
        1958:  q   <=  32'b10111111010110110000011001000010 ;
        1959:  q   <=  32'b00111011111101111010010111110001 ;
        1960:  q   <=  32'b10111111011100000000010110011110 ;
        1961:  q   <=  32'b10111111001011100111101010110010 ;
        1962:  q   <=  32'b10111110100001010011000011111110 ;
        1963:  q   <=  32'b10111110011010100100100101010100 ;
        1964:  q   <=  32'b10111111000001100101101000100100 ;
        1965:  q   <=  32'b00111111100100000110110010111101 ;
        1966:  q   <=  32'b00111111000011001101010111101101 ;
        1967:  q   <=  32'b00111111111011010111010101110111 ;
        1968:  q   <=  32'b10111110100011011111101000011011 ;
        1969:  q   <=  32'b00111111100010001000011101011011 ;
        1970:  q   <=  32'b11000000000001100101100111101101 ;
        1971:  q   <=  32'b00111111001000110111001110101100 ;
        1972:  q   <=  32'b00111110101111100011000010111000 ;
        1973:  q   <=  32'b10111110101111111001010001101101 ;
        1974:  q   <=  32'b00111111001100100000001001011001 ;
        1975:  q   <=  32'b00111111011000001010110001000110 ;
        1976:  q   <=  32'b00111111100001000100110100110000 ;
        1977:  q   <=  32'b00111110110101101110111011100011 ;
        1978:  q   <=  32'b00111111000110011101111110101100 ;
        1979:  q   <=  32'b10111111001011001000110001110110 ;
        1980:  q   <=  32'b10111111100011000010111011001110 ;
        1981:  q   <=  32'b10111110100010010000010100001111 ;
        1982:  q   <=  32'b00111110001111110000011100001111 ;
        1983:  q   <=  32'b00111111011100110111000100011100 ;
        1984:  q   <=  32'b10111111010010100101111101101111 ;
        1985:  q   <=  32'b10111110111110101001110011011011 ;
        1986:  q   <=  32'b01000000001111100101110111000111 ;
        1987:  q   <=  32'b10111111000111110110000111000001 ;
        1988:  q   <=  32'b00111111111101011100110001111101 ;
        1989:  q   <=  32'b00111111011101100000110111011011 ;
        1990:  q   <=  32'b10111111000011101100110000110000 ;
        1991:  q   <=  32'b10111101110110100011100110010110 ;
        1992:  q   <=  32'b10111110010111000101001100111010 ;
        1993:  q   <=  32'b00111110111100100110110100111101 ;
        1994:  q   <=  32'b00111111101011101100110101010010 ;
        1995:  q   <=  32'b10111111110100011010001110001101 ;
        1996:  q   <=  32'b01000000000000011000010011000110 ;
        1997:  q   <=  32'b00111111010001110001110100110010 ;
        1998:  q   <=  32'b10111111000011001000010011010110 ;
        1999:  q   <=  32'b10111110000000010000100100011111 ;
        2000:  q   <=  32'b00111110100110010110001010011010 ;
        2001:  q   <=  32'b00111110100101111010001110111111 ;
        2002:  q   <=  32'b00111111100110011011001101000001 ;
        2003:  q   <=  32'b00111111100010111000101011001000 ;
        2004:  q   <=  32'b10111110101101111010011111110010 ;
        2005:  q   <=  32'b10111110000001010000101110111111 ;
        2006:  q   <=  32'b00111111001110111101011000111000 ;
        2007:  q   <=  32'b00111101111101100111000001100101 ;
        2008:  q   <=  32'b00111111100100010111001101001101 ;
        2009:  q   <=  32'b10111111001011111101000001011100 ;
        2010:  q   <=  32'b00111110111100011000000001101010 ;
        2011:  q   <=  32'b00111110100100111010000110011111 ;
        2012:  q   <=  32'b00111111101100100010100001001100 ;
        2013:  q   <=  32'b10111111101011000011100101101000 ;
        2014:  q   <=  32'b00111010010000111110110110010100 ;
        2015:  q   <=  32'b00111101010110110001110101011111 ;
        2016:  q   <=  32'b11000000000101011110000111000110 ;
        2017:  q   <=  32'b00111111100111111100000110010100 ;
        2018:  q   <=  32'b01000000001100111100101001110100 ;
        2019:  q   <=  32'b10111110011011011100000111011110 ;
        2020:  q   <=  32'b00111110100100101111010111100000 ;
        2021:  q   <=  32'b10111110111011011110000010100011 ;
        2022:  q   <=  32'b00111110110001001100010101001100 ;
        2023:  q   <=  32'b10111110110000100111100011000000 ;
        2024:  q   <=  32'b10111101110100000111000100011010 ;
        2025:  q   <=  32'b00111111110011110001111110010011 ;
        2026:  q   <=  32'b10111111010110001110010000001110 ;
        2027:  q   <=  32'b10111111000100110110110100010100 ;
        2028:  q   <=  32'b10111101100110110111100001010111 ;
        2029:  q   <=  32'b10111110000001111010011010100010 ;
        2030:  q   <=  32'b00111111101110000011101101001100 ;
        2031:  q   <=  32'b01000000000000100000000000110110 ;
        2032:  q   <=  32'b10111111011110100110101101101011 ;
        2033:  q   <=  32'b10111111001001000001101000100000 ;
        2034:  q   <=  32'b00111111000001010011110111100100 ;
        2035:  q   <=  32'b10111110110000101110101100011100 ;
        2036:  q   <=  32'b00111111111111110001010111000101 ;
        2037:  q   <=  32'b00111111110100010110010000110010 ;
        2038:  q   <=  32'b00111111000011110001101111011100 ;
        2039:  q   <=  32'b00111111000100000100101010001101 ;
        2040:  q   <=  32'b10111110101011010100001001010010 ;
        2041:  q   <=  32'b00111111010000110111111001100100 ;
        2042:  q   <=  32'b00111111100100000101000000000111 ;
        2043:  q   <=  32'b00111110000100001111100000001000 ;
        2044:  q   <=  32'b00111111111101101100110100011001 ;
        2045:  q   <=  32'b00111111001010111010111011101101 ;
        2046:  q   <=  32'b10111101111000011000001000000000 ;
        2047:  q   <=  32'b00111110101111011110111011000011 ;
        2048:  q   <=  32'b00111111100011000101110100110111 ;
        2049:  q   <=  32'b10111110110010111101110000001000 ;
        2050:  q   <=  32'b10111101101011110000011011111101 ;
        2051:  q   <=  32'b01000000000101111110001111110000 ;
        2052:  q   <=  32'b10111110111100101010010111000110 ;
        2053:  q   <=  32'b00111111011100100100001101100100 ;
        2054:  q   <=  32'b00111111010100010111001100001001 ;
        2055:  q   <=  32'b00111111110010110110001101100101 ;
        2056:  q   <=  32'b00111111000001101010100010111000 ;
        2057:  q   <=  32'b11000000000111011100010111001011 ;
        2058:  q   <=  32'b10111111010110100011111101000101 ;
        2059:  q   <=  32'b00111111000000110000000100010111 ;
        2060:  q   <=  32'b00111110100000111111101100010010 ;
        2061:  q   <=  32'b00111111111110110011000101111001 ;
        2062:  q   <=  32'b00111111101101000000001000100000 ;
        2063:  q   <=  32'b00111110111111100110000011111101 ;
        2064:  q   <=  32'b00111101101010011010001100010001 ;
        2065:  q   <=  32'b10111111110001100011010010000101 ;
        2066:  q   <=  32'b00111111111011100111110000000011 ;
        2067:  q   <=  32'b00111110000010010011111001000110 ;
        2068:  q   <=  32'b10111111110001011110001101101001 ;
        2069:  q   <=  32'b00111110110111011101011100110000 ;
        2070:  q   <=  32'b00111101110100101101100110101001 ;
        2071:  q   <=  32'b10111111000100100000001000110011 ;
        2072:  q   <=  32'b00111110111111000111001010100100 ;
        2073:  q   <=  32'b10111111001101010001111110010110 ;
        2074:  q   <=  32'b10111111101011001000110000010101 ;
        2075:  q   <=  32'b10111111111000001000110011110011 ;
        2076:  q   <=  32'b10111110101110100100010100101010 ;
        2077:  q   <=  32'b10111111001000001000100100111011 ;
        2078:  q   <=  32'b00111110111000010101101101011111 ;
        2079:  q   <=  32'b10111111110000000101011010001011 ;
        2080:  q   <=  32'b10111110010101010011101110101100 ;
        2081:  q   <=  32'b10111111110000001010011111110011 ;
        2082:  q   <=  32'b00111111111001111010010110010110 ;
        2083:  q   <=  32'b10111101111011111000111101010000 ;
        2084:  q   <=  32'b00111111100111001111010001101010 ;
        2085:  q   <=  32'b00111110111111010110100100110000 ;
        2086:  q   <=  32'b00111111011010001001100110101100 ;
        2087:  q   <=  32'b10111111100100111011110101110001 ;
        2088:  q   <=  32'b00111111101000001111011110010100 ;
        2089:  q   <=  32'b00111111101110011110110010010101 ;
        2090:  q   <=  32'b11000000000001001110101001111010 ;
        2091:  q   <=  32'b10111110001101001011100101000101 ;
        2092:  q   <=  32'b10111111001001101110111011011011 ;
        2093:  q   <=  32'b00111110001000000100101001100101 ;
        2094:  q   <=  32'b10111111010110011010100001100101 ;
        2095:  q   <=  32'b00111110100011101101111100011011 ;
        2096:  q   <=  32'b00111111000110001101101100100010 ;
        2097:  q   <=  32'b00111110011110101001011100000100 ;
        2098:  q   <=  32'b10111101111100100101111110100111 ;
        2099:  q   <=  32'b10111111101001010000101101010001 ;
        2100:  q   <=  32'b00111101011010111100011111011010 ;
        2101:  q   <=  32'b10111111000001010101101111011011 ;
        2102:  q   <=  32'b10111111101000111011011100100111 ;
        2103:  q   <=  32'b10111101011001100100111010000110 ;
        2104:  q   <=  32'b10111110010101101011011001101101 ;
        2105:  q   <=  32'b00111110010001001011011001000101 ;
        2106:  q   <=  32'b00111111011111100000100101111101 ;
        2107:  q   <=  32'b00111111000100111000010010111101 ;
        2108:  q   <=  32'b00111111101001110010001111101100 ;
        2109:  q   <=  32'b10111111001110101011001111001001 ;
        2110:  q   <=  32'b10111111010111010101010011000100 ;
        2111:  q   <=  32'b10111101110000100110010111101111 ;
        2112:  q   <=  32'b00111111101100010000110100100111 ;
        2113:  q   <=  32'b00111111101001101101111100000111 ;
        2114:  q   <=  32'b10111110000000001101010011101000 ;
        2115:  q   <=  32'b10111111000110001100110010111000 ;
        2116:  q   <=  32'b10111111110000101010010010001001 ;
        2117:  q   <=  32'b00111111001010111111110111001111 ;
        2118:  q   <=  32'b00111100101110110010001111110010 ;
        2119:  q   <=  32'b10111111100101101100000111000110 ;
        2120:  q   <=  32'b10111110101010110100110111010100 ;
        2121:  q   <=  32'b10111111111010100010101110010110 ;
        2122:  q   <=  32'b00111110110111000010011110011000 ;
        2123:  q   <=  32'b10111110001100100010101101010111 ;
        2124:  q   <=  32'b00111111110100001100110010001101 ;
        2125:  q   <=  32'b10111111101011100000000110111100 ;
        2126:  q   <=  32'b00111111011110000111001100100000 ;
        2127:  q   <=  32'b00111110000100110001011001010000 ;
        2128:  q   <=  32'b00111101101010010010110000010010 ;
        2129:  q   <=  32'b00111111001101110111011101001010 ;
        2130:  q   <=  32'b00111111100110001100010000010100 ;
        2131:  q   <=  32'b10111111100010010001100010001110 ;
        2132:  q   <=  32'b00111111101010001101000111001001 ;
        2133:  q   <=  32'b10111111100110101110000101100010 ;
        2134:  q   <=  32'b10111111100010010111110010011000 ;
        2135:  q   <=  32'b10111111001011000010110011100101 ;
        2136:  q   <=  32'b00111111001111001000100011001001 ;
        2137:  q   <=  32'b10111111100010001111010001111000 ;
        2138:  q   <=  32'b00111110101010110101111111000111 ;
        2139:  q   <=  32'b00111110110100101110001001000110 ;
        2140:  q   <=  32'b00111110000111011101000110101110 ;
        2141:  q   <=  32'b00111111000011011111100001011000 ;
        2142:  q   <=  32'b10111111100101100001111111001110 ;
        2143:  q   <=  32'b00111111100000001111100010011001 ;
        2144:  q   <=  32'b00111101111010000111110101010010 ;
        2145:  q   <=  32'b00111111001110101110010010011101 ;
        2146:  q   <=  32'b10111111011110111100011101101101 ;
        2147:  q   <=  32'b00111101010101010001111100001010 ;
        2148:  q   <=  32'b00111111011000001010101001011010 ;
        2149:  q   <=  32'b00111111100000011100111101011111 ;
        2150:  q   <=  32'b10111101101011001011111011011100 ;
        2151:  q   <=  32'b10111111111011010100000010000101 ;
        2152:  q   <=  32'b10111111100011000110010010011110 ;
        2153:  q   <=  32'b00111110010111111101111111101011 ;
        2154:  q   <=  32'b00111111010010110101001110110010 ;
        2155:  q   <=  32'b00111110111011010001111010011101 ;
        2156:  q   <=  32'b10111111000111001101010101010010 ;
        2157:  q   <=  32'b01000000000011111010010000111111 ;
        2158:  q   <=  32'b00111101100101000010101011111011 ;
        2159:  q   <=  32'b00111111010111011001001001011001 ;
        2160:  q   <=  32'b10111110110101001101011000101010 ;
        2161:  q   <=  32'b10111111100011101011011001001010 ;
        2162:  q   <=  32'b00111111001011110110110010110011 ;
        2163:  q   <=  32'b00111111100001001101001001111001 ;
        2164:  q   <=  32'b00111111111010010011111000111010 ;
        2165:  q   <=  32'b10111111000001110110101111001010 ;
        2166:  q   <=  32'b10111111110100000110000100110110 ;
        2167:  q   <=  32'b00111111110011110000001111000100 ;
        2168:  q   <=  32'b00111110100001110011110011101110 ;
        2169:  q   <=  32'b10111111100100000100011001010011 ;
        2170:  q   <=  32'b10111111000011110010011000100110 ;
        2171:  q   <=  32'b10111111010011110001000001111001 ;
        2172:  q   <=  32'b00111111100101001001101111001001 ;
        2173:  q   <=  32'b00111111000101111001010000110101 ;
        2174:  q   <=  32'b00111110011110001001001011011000 ;
        2175:  q   <=  32'b00111110011101100011111110111010 ;
        2176:  q   <=  32'b10111111010100100100110111011001 ;
        2177:  q   <=  32'b00111111011111100011110010011000 ;
        2178:  q   <=  32'b00111110101100010101101010100110 ;
        2179:  q   <=  32'b10111110100001011011001101001011 ;
        2180:  q   <=  32'b10111110001111010010010101100001 ;
        2181:  q   <=  32'b10111101110100000101101001110000 ;
        2182:  q   <=  32'b10111111011000110001010101000010 ;
        2183:  q   <=  32'b00111111001111011100101011100011 ;
        2184:  q   <=  32'b00111111101100100011001111011110 ;
        2185:  q   <=  32'b01000000000111100101010001100001 ;
        2186:  q   <=  32'b00111111000000010000000011011001 ;
        2187:  q   <=  32'b10111111010100101000111000010101 ;
        2188:  q   <=  32'b00111110010011011100111000110001 ;
        2189:  q   <=  32'b10111111100000001110011100011000 ;
        2190:  q   <=  32'b10111111000111001111100011001111 ;
        2191:  q   <=  32'b10111111001010001011000111010011 ;
        2192:  q   <=  32'b10111111010101010100111010000100 ;
        2193:  q   <=  32'b00111110110000011010000010110111 ;
        2194:  q   <=  32'b10111111100011101100001110001011 ;
        2195:  q   <=  32'b00111111001010101101000001010100 ;
        2196:  q   <=  32'b00111111010010111001101011101110 ;
        2197:  q   <=  32'b00111111100001001100110010001000 ;
        2198:  q   <=  32'b10111100101001110101111101010001 ;
        2199:  q   <=  32'b00111111000111100111001110110101 ;
        2200:  q   <=  32'b00111111111001101100101011001000 ;
        2201:  q   <=  32'b00111101010110010000111110000011 ;
        2202:  q   <=  32'b10111110001101100010100011010001 ;
        2203:  q   <=  32'b00111111111000101110000010110101 ;
        2204:  q   <=  32'b11000000001000001001000000111101 ;
        2205:  q   <=  32'b10111110111010011100011000001110 ;
        2206:  q   <=  32'b01000000000110111000101101001110 ;
        2207:  q   <=  32'b10111110111100010110001001101110 ;
        2208:  q   <=  32'b10111111000011110111000110110000 ;
        2209:  q   <=  32'b10111111100111001111110011100010 ;
        2210:  q   <=  32'b00111111010010101111111011001011 ;
        2211:  q   <=  32'b11000000000001110000100101000011 ;
        2212:  q   <=  32'b10111111010011001010010100101000 ;
        2213:  q   <=  32'b00111111000100010010010101000111 ;
        2214:  q   <=  32'b10111010101111010001111110100110 ;
        2215:  q   <=  32'b00111111000111111011100110000110 ;
        2216:  q   <=  32'b00111110000000010111100110110100 ;
        2217:  q   <=  32'b00111111001011100100110101011010 ;
        2218:  q   <=  32'b10111111101001001100101000001011 ;
        2219:  q   <=  32'b00111110010111110101000110100010 ;
        2220:  q   <=  32'b10111111110010001000010101000101 ;
        2221:  q   <=  32'b00111111010010001000010100101010 ;
        2222:  q   <=  32'b10111110100111110000001100000100 ;
        2223:  q   <=  32'b00111111001001111100001101010111 ;
        2224:  q   <=  32'b10111111000010011001011101110101 ;
        2225:  q   <=  32'b00111110101010000100001111110010 ;
        2226:  q   <=  32'b00111111100001101110101111010100 ;
        2227:  q   <=  32'b10111111111111010110011011001001 ;
        2228:  q   <=  32'b10111111111011110000011010010011 ;
        2229:  q   <=  32'b10111111111010101000101010100001 ;
        2230:  q   <=  32'b00111111010110010011110101010101 ;
        2231:  q   <=  32'b00111110110011110111010010110100 ;
        2232:  q   <=  32'b10111111001100111101010000101000 ;
        2233:  q   <=  32'b00111111101111111110000010111101 ;
        2234:  q   <=  32'b00111110000011010001101000011000 ;
        2235:  q   <=  32'b10111111110010110001110011110110 ;
        2236:  q   <=  32'b10111111100000100111001101011100 ;
        2237:  q   <=  32'b10111111101100010100111101010110 ;
        2238:  q   <=  32'b00111111011101000111001101101111 ;
        2239:  q   <=  32'b10111111000110011110001100000101 ;
        2240:  q   <=  32'b10111111100101100000000010000100 ;
        2241:  q   <=  32'b10111111000100111011110110000000 ;
        2242:  q   <=  32'b10111111010101100010000001001111 ;
        2243:  q   <=  32'b00111111010110100101110000110110 ;
        2244:  q   <=  32'b00111110111101000110010011000000 ;
        2245:  q   <=  32'b00111110100110101100100110110010 ;
        2246:  q   <=  32'b00111110110101001110000010011101 ;
        2247:  q   <=  32'b00111101001100000000011001011111 ;
        2248:  q   <=  32'b10111111011100101110100000001011 ;
        2249:  q   <=  32'b00111111000010101010011011011000 ;
        2250:  q   <=  32'b10111111010100100011010101110110 ;
        2251:  q   <=  32'b10111111100010010011010000101111 ;
        2252:  q   <=  32'b10111111100010010111101111010101 ;
        2253:  q   <=  32'b00111111010111101001101100000011 ;
        2254:  q   <=  32'b00111111011110110010011000101111 ;
        2255:  q   <=  32'b10111111111000010010000100110000 ;
        2256:  q   <=  32'b10111110000101111010011001110111 ;
        2257:  q   <=  32'b00111110100000001111111010000010 ;
        2258:  q   <=  32'b10111111000111000100001000101010 ;
        2259:  q   <=  32'b00111111010000101100111110010010 ;
        2260:  q   <=  32'b00111110100000100100010010010101 ;
        2261:  q   <=  32'b10111110000111001000000001101110 ;
        2262:  q   <=  32'b10111111000011101011001001111010 ;
        2263:  q   <=  32'b00111111001011010101000100000111 ;
        2264:  q   <=  32'b00111111010110010110101110001110 ;
        2265:  q   <=  32'b00111110111100000100100100000111 ;
        2266:  q   <=  32'b10111110011101011000100101010101 ;
        2267:  q   <=  32'b00111111011010111100010110110011 ;
        2268:  q   <=  32'b10111111011010000010100101100000 ;
        2269:  q   <=  32'b00111110000100111110100000111101 ;
        2270:  q   <=  32'b00111111101100101011110110000111 ;
        2271:  q   <=  32'b10111110010000100100000001100100 ;
        2272:  q   <=  32'b10111111010110000000010110100001 ;
        2273:  q   <=  32'b00111111111110001100001010010011 ;
        2274:  q   <=  32'b10111110011111001101100100000000 ;
        2275:  q   <=  32'b00111110111000100001101111100111 ;
        2276:  q   <=  32'b10111111010011011011100101111011 ;
        2277:  q   <=  32'b00111110100100110100000110001011 ;
        2278:  q   <=  32'b00111110111011110001110011111110 ;
        2279:  q   <=  32'b00111011100101010111100110001101 ;
        2280:  q   <=  32'b00111110101001101111010101010000 ;
        2281:  q   <=  32'b00111111100110100010111111100101 ;
        2282:  q   <=  32'b10111111101100111011101000010001 ;
        2283:  q   <=  32'b00111110010100100111111101000000 ;
        2284:  q   <=  32'b10111111111111101101111110000000 ;
        2285:  q   <=  32'b00111100111010001011100111011010 ;
        2286:  q   <=  32'b00111111111101110001101100100001 ;
        2287:  q   <=  32'b00111111011100001110111001010111 ;
        2288:  q   <=  32'b10111011111000101110011010000001 ;
        2289:  q   <=  32'b10111110101011010010111000000010 ;
        2290:  q   <=  32'b00111111000001110011110001101101 ;
        2291:  q   <=  32'b00111111100001110100100001111100 ;
        2292:  q   <=  32'b00111100011100011000001010100000 ;
        2293:  q   <=  32'b00111111110011101011000001111111 ;
        2294:  q   <=  32'b10111111010100001101101111011110 ;
        2295:  q   <=  32'b10111111111111111011011010010010 ;
        2296:  q   <=  32'b10111111001111111000100101111000 ;
        2297:  q   <=  32'b10111110010011000001011001011010 ;
        2298:  q   <=  32'b10111110101111101101101001101000 ;
        2299:  q   <=  32'b10111111010110001110110101010000 ;
        2300:  q   <=  32'b00111111101010110010101010011101 ;
        2301:  q   <=  32'b10111111110011101110001101111011 ;
        2302:  q   <=  32'b10111110111110111100111110000100 ;
        2303:  q   <=  32'b10111111011110000010010000100101 ;
        2304:  q   <=  32'b10111110111100101011111001000101 ;
        2305:  q   <=  32'b10111111001010101000100110110110 ;
        2306:  q   <=  32'b00111110111101001110110110000110 ;
        2307:  q   <=  32'b10111111100001010100000101100100 ;
        2308:  q   <=  32'b10111111010100100001011010110110 ;
        2309:  q   <=  32'b00111101110011110001110100001001 ;
        2310:  q   <=  32'b00111111100010101011111111110000 ;
        2311:  q   <=  32'b10111111111011010110000100100110 ;
        2312:  q   <=  32'b00111111111001100101111001001100 ;
        2313:  q   <=  32'b10111111011000001101110100100011 ;
        2314:  q   <=  32'b00111111001001011101000111001111 ;
        2315:  q   <=  32'b00111111100001100101100000100101 ;
        2316:  q   <=  32'b00111111101010010101101100011111 ;
        2317:  q   <=  32'b10111111000001000111000110100011 ;
        2318:  q   <=  32'b00111100110001110011000000100101 ;
        2319:  q   <=  32'b10111110001001100100001110000000 ;
        2320:  q   <=  32'b10111111000110110000110010011010 ;
        2321:  q   <=  32'b00111110100010110001110110001010 ;
        2322:  q   <=  32'b00111110101101111010000000011011 ;
        2323:  q   <=  32'b10111110101101000110001010100101 ;
        2324:  q   <=  32'b00111110000001111000100101011100 ;
        2325:  q   <=  32'b01000000001010110001101111110110 ;
        2326:  q   <=  32'b10111011111101111110110011010111 ;
        2327:  q   <=  32'b00111111001101011101011001101001 ;
        2328:  q   <=  32'b10111110111011001101000111110101 ;
        2329:  q   <=  32'b10111111000001110010001100000001 ;
        2330:  q   <=  32'b10111110101100010000101100000000 ;
        2331:  q   <=  32'b00111111000100001000011011011011 ;
        2332:  q   <=  32'b10111111010011010011000110101011 ;
        2333:  q   <=  32'b10111111111011010010110101011100 ;
        2334:  q   <=  32'b00111101010110011111100100001001 ;
        2335:  q   <=  32'b10111110110111110111000111010000 ;
        2336:  q   <=  32'b00111110100011110101110100100011 ;
        2337:  q   <=  32'b00111101101011010100010111011001 ;
        2338:  q   <=  32'b00111111001110101010011110001011 ;
        2339:  q   <=  32'b00111111011001101001011111000001 ;
        2340:  q   <=  32'b10111111101010011010111010000100 ;
        2341:  q   <=  32'b10111111110000110010010101100110 ;
        2342:  q   <=  32'b00111111000000001001111101111000 ;
        2343:  q   <=  32'b00111110100111001101111101010110 ;
        2344:  q   <=  32'b10111111011100000110110011010001 ;
        2345:  q   <=  32'b00111111100111100110001100110001 ;
        2346:  q   <=  32'b00111101000001110011011110000000 ;
        2347:  q   <=  32'b00111101111111010001000101100010 ;
        2348:  q   <=  32'b00111110100011000100000111001000 ;
        2349:  q   <=  32'b00111111010000010001000100000010 ;
        2350:  q   <=  32'b00111111110000110010001010111011 ;
        2351:  q   <=  32'b10111110100001100010000110101111 ;
        2352:  q   <=  32'b10111111110111011000011100001001 ;
        2353:  q   <=  32'b00111111100000011011100100110010 ;
        2354:  q   <=  32'b10111111011011011000000000011100 ;
        2355:  q   <=  32'b00111111100111110011000011101010 ;
        2356:  q   <=  32'b10111111000101101110100010111011 ;
        2357:  q   <=  32'b00111111101111101110100011011111 ;
        2358:  q   <=  32'b10111111010011100101010010010100 ;
        2359:  q   <=  32'b10111111100011100110100110100101 ;
        2360:  q   <=  32'b00111111011101001111100111111101 ;
        2361:  q   <=  32'b10111111101011100111100001111001 ;
        2362:  q   <=  32'b00111111001011100011101011010000 ;
        2363:  q   <=  32'b00111110111000000010101001101010 ;
        2364:  q   <=  32'b10111110000100101011010010111010 ;
        2365:  q   <=  32'b10111110101011101101110101011001 ;
        2366:  q   <=  32'b01000000000000111011001100101011 ;
        2367:  q   <=  32'b10111110101111111100001100001110 ;
        2368:  q   <=  32'b10111110010000101100010010100000 ;
        2369:  q   <=  32'b10111111011100000101000011000100 ;
        2370:  q   <=  32'b10111111010100000011111100010001 ;
        2371:  q   <=  32'b10111111000101010110100000001001 ;
        2372:  q   <=  32'b00111111110110101101000110111010 ;
        2373:  q   <=  32'b10111110110001111110010100011011 ;
        2374:  q   <=  32'b10111111001100001010100000011111 ;
        2375:  q   <=  32'b10111110111001010111110100101111 ;
        2376:  q   <=  32'b00111111001101101110000101011110 ;
        2377:  q   <=  32'b10111111101010000110100111100001 ;
        2378:  q   <=  32'b00111111001000001000101100010010 ;
        2379:  q   <=  32'b10111111101010100110011111011110 ;
        2380:  q   <=  32'b10111110000001011111110100001110 ;
        2381:  q   <=  32'b10111111111010011101011110111011 ;
        2382:  q   <=  32'b00111111000010010011001000110110 ;
        2383:  q   <=  32'b00111111001100010101111110010100 ;
        2384:  q   <=  32'b10111111001100000000001101000010 ;
        2385:  q   <=  32'b00111110101000101001100101001010 ;
        2386:  q   <=  32'b00111110001001101100000000100100 ;
        2387:  q   <=  32'b00111111100101000101110111101000 ;
        2388:  q   <=  32'b00111110000000110111100000101000 ;
        2389:  q   <=  32'b00111111100001010000110011110110 ;
        2390:  q   <=  32'b10111101111011110010010110110101 ;
        2391:  q   <=  32'b10111111001001011111011011001001 ;
        2392:  q   <=  32'b10111101000110111001001000101110 ;
        2393:  q   <=  32'b10111110010011000001101111001110 ;
        2394:  q   <=  32'b00111111011000011011010100011101 ;
        2395:  q   <=  32'b10111101011001011111011101010011 ;
        2396:  q   <=  32'b10111111010101110101101101101110 ;
        2397:  q   <=  32'b10111110000111101000111101100010 ;
        2398:  q   <=  32'b00111111100110000010001111011110 ;
        2399:  q   <=  32'b10111110110101000110111010111010 ;
        2400:  q   <=  32'b10111111001010001001101100011011 ;
        2401:  q   <=  32'b00111111011110111110011011001111 ;
        2402:  q   <=  32'b00111101110011110101000001011100 ;
        2403:  q   <=  32'b10111110101110011011010010010011 ;
        2404:  q   <=  32'b10111111001111010010001111010010 ;
        2405:  q   <=  32'b10111111101111010110101101111001 ;
        2406:  q   <=  32'b00111110000111010000110101111011 ;
        2407:  q   <=  32'b10111110101000100101000000011101 ;
        2408:  q   <=  32'b00111110101000110100100101000000 ;
        2409:  q   <=  32'b10111111101110100111000000011110 ;
        2410:  q   <=  32'b00111111101010010011000111011111 ;
        2411:  q   <=  32'b00111110111110010111001011001011 ;
        2412:  q   <=  32'b10111111110010001000011100110101 ;
        2413:  q   <=  32'b00111111100001110100110110111010 ;
        2414:  q   <=  32'b10111111000101100110101101111111 ;
        2415:  q   <=  32'b00111110100110101011110011001010 ;
        2416:  q   <=  32'b00111110011000001011101010111111 ;
        2417:  q   <=  32'b10111111011000001101000111001001 ;
        2418:  q   <=  32'b11000000001101110010000100101100 ;
        2419:  q   <=  32'b00111111000010010001101000100110 ;
        2420:  q   <=  32'b10111110101011110001111110000011 ;
        2421:  q   <=  32'b10111111000110010000110101000111 ;
        2422:  q   <=  32'b00111110110101100111101110111001 ;
        2423:  q   <=  32'b10111111001100001000111011101010 ;
        2424:  q   <=  32'b00111111001010111101001100101101 ;
        2425:  q   <=  32'b00111110000110101000010011011101 ;
        2426:  q   <=  32'b10111111011111011100011100010011 ;
        2427:  q   <=  32'b00111111010101100011101001111100 ;
        2428:  q   <=  32'b00111110111100101111001011010110 ;
        2429:  q   <=  32'b00111111101000000100011011111000 ;
        2430:  q   <=  32'b10111111011001001000001011101011 ;
        2431:  q   <=  32'b10111111011001010011000010110001 ;
        2432:  q   <=  32'b00111110101000000110110001000001 ;
        2433:  q   <=  32'b00111111001010101100001010101111 ;
        2434:  q   <=  32'b00111111010100111111111101110010 ;
        2435:  q   <=  32'b00111011110101010100101111001000 ;
        2436:  q   <=  32'b10111110011100011000110110111001 ;
        2437:  q   <=  32'b00111111001001110001111101001000 ;
        2438:  q   <=  32'b00111111111110110111010111001101 ;
        2439:  q   <=  32'b00111111011000100111010000011011 ;
        2440:  q   <=  32'b00111101101011010010000110110110 ;
        2441:  q   <=  32'b10111111000100110001001101011010 ;
        2442:  q   <=  32'b00111110111111111101111101010000 ;
        2443:  q   <=  32'b10111110111101111101110010001010 ;
        2444:  q   <=  32'b00111110011101000010101100010111 ;
        2445:  q   <=  32'b00111111010001110011101101000110 ;
        2446:  q   <=  32'b00111111011011001001110100100110 ;
        2447:  q   <=  32'b00111111000101101001000000110100 ;
        2448:  q   <=  32'b00111111101100000110000000100110 ;
        2449:  q   <=  32'b00111111111011001111010001001000 ;
        2450:  q   <=  32'b10111111111100101110011010101101 ;
        2451:  q   <=  32'b10111111111000111010101111101100 ;
        2452:  q   <=  32'b10111111011011000011001000110111 ;
        2453:  q   <=  32'b10111111111111111011110000010011 ;
        2454:  q   <=  32'b10111110101101101101010111010001 ;
        2455:  q   <=  32'b10111110101011000011110010111000 ;
        2456:  q   <=  32'b00111110100000000011011111010110 ;
        2457:  q   <=  32'b00111110100100101000001111010000 ;
        2458:  q   <=  32'b10111111001011111010100010111110 ;
        2459:  q   <=  32'b10111111010100000011010101100000 ;
        2460:  q   <=  32'b00111111010010110001110001101110 ;
        2461:  q   <=  32'b10111110110000111000111001010100 ;
        2462:  q   <=  32'b10111111101011111000001110011110 ;
        2463:  q   <=  32'b00111100001010001110000010011000 ;
        2464:  q   <=  32'b00111110010100010000011111111101 ;
        2465:  q   <=  32'b10111110110100100111000111101111 ;
        2466:  q   <=  32'b00111111001010011101111100100101 ;
        2467:  q   <=  32'b00111110011001110011001101101110 ;
        2468:  q   <=  32'b10111110010110011111001110001011 ;
        2469:  q   <=  32'b10111101001101000101110110011000 ;
        2470:  q   <=  32'b00111110111010101001011011001110 ;
        2471:  q   <=  32'b10111110111000100000000101110101 ;
        2472:  q   <=  32'b10111111100001110000100001111110 ;
        2473:  q   <=  32'b10111110000111110101000101111010 ;
        2474:  q   <=  32'b00111110000001000011111101010110 ;
        2475:  q   <=  32'b00111111000000100110100111100101 ;
        2476:  q   <=  32'b10111100111101101100010110011110 ;
        2477:  q   <=  32'b10111110111010100010101110111101 ;
        2478:  q   <=  32'b00111111000110001010100101110011 ;
        2479:  q   <=  32'b10111101111010001000000110011010 ;
        2480:  q   <=  32'b00111111010011101001100100100110 ;
        2481:  q   <=  32'b10111101101101111110101001111111 ;
        2482:  q   <=  32'b10111011110011100010111000101100 ;
        2483:  q   <=  32'b10111101101111000010000101110010 ;
        2484:  q   <=  32'b10111111011010111101011001000101 ;
        2485:  q   <=  32'b10111111011011010100110010110010 ;
        2486:  q   <=  32'b10111111011101100001001010001110 ;
        2487:  q   <=  32'b00111111111001000111010101001101 ;
        2488:  q   <=  32'b10111110010011001111111001010111 ;
        2489:  q   <=  32'b00111111011100001011111011010001 ;
        2490:  q   <=  32'b00111110101100101100010010011110 ;
        2491:  q   <=  32'b00111111111011011111110011100101 ;
        2492:  q   <=  32'b00111111011011010101010010010110 ;
        2493:  q   <=  32'b10111111100111010000110100100110 ;
        2494:  q   <=  32'b10111110101001111000101111100011 ;
        2495:  q   <=  32'b00111111011001000100001011110000 ;
        2496:  q   <=  32'b00111110100100111000110100001111 ;
        2497:  q   <=  32'b01000000000100001111100011110110 ;
        2498:  q   <=  32'b10111101010001000010100010100110 ;
        2499:  q   <=  32'b10111111110001101010001101111011 ;
        2500:  q   <=  32'b00111110111000110101111011100011 ;
        2501:  q   <=  32'b10111111011010010110110011110110 ;
        2502:  q   <=  32'b00111101010010100111101111111100 ;
        2503:  q   <=  32'b00111111100010011111110101101000 ;
        2504:  q   <=  32'b00111110100111011100100110011011 ;
        2505:  q   <=  32'b00111110100110010110101000111001 ;
        2506:  q   <=  32'b10111110010010011111001110100010 ;
        2507:  q   <=  32'b10111110000101011110111111000011 ;
        2508:  q   <=  32'b10111101110100110001011011010001 ;
        2509:  q   <=  32'b11000000001100110010001010000101 ;
        2510:  q   <=  32'b00111110110010010101101101011101 ;
        2511:  q   <=  32'b00111111011111011000000011010110 ;
        2512:  q   <=  32'b10111111101001100001100011010101 ;
        2513:  q   <=  32'b10111111110000101100111111011011 ;
        2514:  q   <=  32'b00111111000111101111101010011000 ;
        2515:  q   <=  32'b10111111110000001111011010000000 ;
        2516:  q   <=  32'b10111111110101101111011010100110 ;
        2517:  q   <=  32'b00111111010010011111101001011000 ;
        2518:  q   <=  32'b10111111001001110111111100001100 ;
        2519:  q   <=  32'b00111111100111110101100011111011 ;
        2520:  q   <=  32'b10111111101001010110100011101011 ;
        2521:  q   <=  32'b10111111000111010100011000110100 ;
        2522:  q   <=  32'b00111110011101110111111011110011 ;
        2523:  q   <=  32'b00111111000011001010001000100101 ;
        2524:  q   <=  32'b00111110111011110110110111000011 ;
        2525:  q   <=  32'b00111110010001000000110101001101 ;
        2526:  q   <=  32'b10111110011010110101000111111101 ;
        2527:  q   <=  32'b10111111000101000100011110001110 ;
        2528:  q   <=  32'b00111110111101100000000110100000 ;
        2529:  q   <=  32'b10111110110001100000111011101101 ;
        2530:  q   <=  32'b00111110110101111101110111111110 ;
        2531:  q   <=  32'b00111111100010110011100111110010 ;
        2532:  q   <=  32'b11000000000011111111010100001101 ;
        2533:  q   <=  32'b00111111111001101111100100110100 ;
        2534:  q   <=  32'b10111111001000011100111010110101 ;
        2535:  q   <=  32'b00111111101010001000000110110011 ;
        2536:  q   <=  32'b00111111110001101001101010010001 ;
        2537:  q   <=  32'b10111111101111000000010100101110 ;
        2538:  q   <=  32'b00111110001101010010111101010100 ;
        2539:  q   <=  32'b01000000010111011101011100110011 ;
        2540:  q   <=  32'b10111110010110111100011100011011 ;
        2541:  q   <=  32'b00111110111110001111101000000111 ;
        2542:  q   <=  32'b00111110101010010110100111000110 ;
        2543:  q   <=  32'b00111111101000100100101010011101 ;
        2544:  q   <=  32'b00111111100010111001010111111000 ;
        2545:  q   <=  32'b10111111011100100100101010010110 ;
        2546:  q   <=  32'b10111110111000001000001011110101 ;
        2547:  q   <=  32'b00111110101011111011101010011110 ;
        2548:  q   <=  32'b10111101011011110011100001100010 ;
        2549:  q   <=  32'b01000000001000100011110100000110 ;
        2550:  q   <=  32'b00111110111000001001011000100010 ;
        2551:  q   <=  32'b00111110111000000000001001010010 ;
        2552:  q   <=  32'b10111111010101100111000111101111 ;
        2553:  q   <=  32'b10111111101001110101110000111110 ;
        2554:  q   <=  32'b00111111010010110100110011101111 ;
        2555:  q   <=  32'b10111110010010011111111110000100 ;
        2556:  q   <=  32'b00111111001001100010111011100001 ;
        2557:  q   <=  32'b10111111010101001101101101111111 ;
        2558:  q   <=  32'b00111111011001010101110100111110 ;
        2559:  q   <=  32'b10111111111010000010000001010010 ;
        2560:  q   <=  32'b00111111110010001000100100010101 ;
        2561:  q   <=  32'b00111111010110001011010001000100 ;
        2562:  q   <=  32'b00111101111000011001100011011011 ;
        2563:  q   <=  32'b10111111100101001001111011111001 ;
        2564:  q   <=  32'b10111110110010111000100111001100 ;
        2565:  q   <=  32'b00111110100000100011001011011101 ;
        2566:  q   <=  32'b00111111100110101001100011011000 ;
        2567:  q   <=  32'b10111111100001000100101100010111 ;
        2568:  q   <=  32'b00111111101001011100011101011110 ;
        2569:  q   <=  32'b01000000001100010010100011101101 ;
        2570:  q   <=  32'b10111110111111011001111000100100 ;
        2571:  q   <=  32'b00111110111100000000001000001000 ;
        2572:  q   <=  32'b10111111001010000100010010011011 ;
        2573:  q   <=  32'b10111111110110111100010101000001 ;
        2574:  q   <=  32'b00111111101111000011100111111000 ;
        2575:  q   <=  32'b00111111001100011011001011111010 ;
        2576:  q   <=  32'b10111111000000101011110100001001 ;
        2577:  q   <=  32'b00111101111010000011011110100100 ;
        2578:  q   <=  32'b10111110011010110101001010010000 ;
        2579:  q   <=  32'b10111111101110110001101000001111 ;
        2580:  q   <=  32'b11000000001110000111100000110010 ;
        2581:  q   <=  32'b10111101010000100110110101100100 ;
        2582:  q   <=  32'b10111110111011001100100001010110 ;
        2583:  q   <=  32'b10111111000100111001111100010000 ;
        2584:  q   <=  32'b10111111010110001001000101100001 ;
        2585:  q   <=  32'b10111111111010001001101100101100 ;
        2586:  q   <=  32'b10111111000001011001000000100011 ;
        2587:  q   <=  32'b00111110001001010100111101110010 ;
        2588:  q   <=  32'b10111111100001111110100101101011 ;
        2589:  q   <=  32'b00111110111001101010011100011101 ;
        2590:  q   <=  32'b10111110100010111010110000110000 ;
        2591:  q   <=  32'b10111101110011111100011101001100 ;
        2592:  q   <=  32'b10111111101101101110110011110001 ;
        2593:  q   <=  32'b10111111010000111011000001010110 ;
        2594:  q   <=  32'b00111110110100011111110110001100 ;
        2595:  q   <=  32'b10111111010010100011100100001000 ;
        2596:  q   <=  32'b00111110001001011000010000110100 ;
        2597:  q   <=  32'b00111111111111010010101111110101 ;
        2598:  q   <=  32'b00111111010010111001011010010100 ;
        2599:  q   <=  32'b00111111100001001100100001101110 ;
        2600:  q   <=  32'b01000000000101110000111110100101 ;
        2601:  q   <=  32'b00111111100101100111001101011000 ;
        2602:  q   <=  32'b00111110110010111010010010100010 ;
        2603:  q   <=  32'b00111111111110011100001010000100 ;
        2604:  q   <=  32'b10111111011001111001011110001111 ;
        2605:  q   <=  32'b10111111001011101010000110000110 ;
        2606:  q   <=  32'b01000000000000010010101110110000 ;
        2607:  q   <=  32'b00111110111010001001111110101011 ;
        2608:  q   <=  32'b10111101001011000111010101101110 ;
        2609:  q   <=  32'b00111110111010101001010011100111 ;
        2610:  q   <=  32'b10111110100001110011110111100110 ;
        2611:  q   <=  32'b10111110100101010111111100010011 ;
        2612:  q   <=  32'b10111110110001100000101001101000 ;
        2613:  q   <=  32'b10111111000011011101001001111011 ;
        2614:  q   <=  32'b10111111011100011001100000100111 ;
        2615:  q   <=  32'b10111101011101010010001101011110 ;
        2616:  q   <=  32'b10111111000100110001111010001010 ;
        2617:  q   <=  32'b00111111101110001000111010110110 ;
        2618:  q   <=  32'b00111110011100010010110111101011 ;
        2619:  q   <=  32'b00111111100000101011110001110111 ;
        2620:  q   <=  32'b10111110000011110010111110111100 ;
        2621:  q   <=  32'b10111101101001110000010001000011 ;
        2622:  q   <=  32'b00111111101000010000111000111010 ;
        2623:  q   <=  32'b00111111101110111111100011101100 ;
        2624:  q   <=  32'b00111101000001101110110011111101 ;
        2625:  q   <=  32'b00111111110110001010001100011111 ;
        2626:  q   <=  32'b00111110111100111001001010110001 ;
        2627:  q   <=  32'b00111110101111001010111111111110 ;
        2628:  q   <=  32'b01000000000011000100100110111101 ;
        2629:  q   <=  32'b00111111110001001001000101010100 ;
        2630:  q   <=  32'b00111111011010000100001000110100 ;
        2631:  q   <=  32'b00111110110011011111010011110111 ;
        2632:  q   <=  32'b10111111000010011101001101100111 ;
        2633:  q   <=  32'b10111101111010111111011000011001 ;
        2634:  q   <=  32'b00111111111010010011011101001100 ;
        2635:  q   <=  32'b11000000000000010110000001011101 ;
        2636:  q   <=  32'b10111111001000110001000011110100 ;
        2637:  q   <=  32'b10111110010000010101010110100001 ;
        2638:  q   <=  32'b00111110000101111101010101101001 ;
        2639:  q   <=  32'b10111111111001000101011000101110 ;
        2640:  q   <=  32'b00111111000001110111000011111000 ;
        2641:  q   <=  32'b00111111001110101100111110110101 ;
        2642:  q   <=  32'b10111111011100001010110010101110 ;
        2643:  q   <=  32'b10111110100001001100000101000010 ;
        2644:  q   <=  32'b10111111100110110101010101101111 ;
        2645:  q   <=  32'b00111111110011111111000100111110 ;
        2646:  q   <=  32'b00111110101111110011110100000100 ;
        2647:  q   <=  32'b10111110100000000111010011100011 ;
        2648:  q   <=  32'b10111111011011001110101010101101 ;
        2649:  q   <=  32'b00111101110010100000111001101101 ;
        2650:  q   <=  32'b00111111110101111001011001111011 ;
        2651:  q   <=  32'b00111110100011001110111011001100 ;
        2652:  q   <=  32'b00111110101101001110001001011000 ;
        2653:  q   <=  32'b10111111100110011010010111101000 ;
        2654:  q   <=  32'b00111110001010100001110110100010 ;
        2655:  q   <=  32'b00111111010001101011001010001001 ;
        2656:  q   <=  32'b10111111101100001101001011100000 ;
        2657:  q   <=  32'b00111111100100000110101101110010 ;
        2658:  q   <=  32'b01000000000111011100100111000011 ;
        2659:  q   <=  32'b10111111110001110110100111010100 ;
        2660:  q   <=  32'b11000000000001000100001111110101 ;
        2661:  q   <=  32'b10111101100101001010111010011011 ;
        2662:  q   <=  32'b00111111010000100101010100100000 ;
        2663:  q   <=  32'b10111101101001110011111110001000 ;
        2664:  q   <=  32'b10111110001000100100011011010010 ;
        2665:  q   <=  32'b00111011110101001110110101111011 ;
        2666:  q   <=  32'b10111111100010000100010100010001 ;
        2667:  q   <=  32'b10111111110100100110101111001111 ;
        2668:  q   <=  32'b00111111110010100111000000111001 ;
        2669:  q   <=  32'b00111110100101011101000110000101 ;
        2670:  q   <=  32'b10111111100110000000001110001110 ;
        2671:  q   <=  32'b00111111100010011011100001001011 ;
        2672:  q   <=  32'b10111111101001100001000001000101 ;
        2673:  q   <=  32'b10111101111110010110001010101011 ;
        2674:  q   <=  32'b00111111001111011010001100110100 ;
        2675:  q   <=  32'b10111111010101110011100101000101 ;
        2676:  q   <=  32'b10111110101100101110110111010110 ;
        2677:  q   <=  32'b00111100111100101011111010110111 ;
        2678:  q   <=  32'b00111111111110011110011101011111 ;
        2679:  q   <=  32'b00111110111010110000010100100001 ;
        2680:  q   <=  32'b10111110110011000111001010011101 ;
        2681:  q   <=  32'b10111110011001101100101100111011 ;
        2682:  q   <=  32'b10111110100011111000000100111110 ;
        2683:  q   <=  32'b00111111101001110100001011000000 ;
        2684:  q   <=  32'b10111110100100011001100110011110 ;
        2685:  q   <=  32'b10111111010010101010110110001001 ;
        2686:  q   <=  32'b00111110011101100110010011001100 ;
        2687:  q   <=  32'b10111101110000011101010111000000 ;
        2688:  q   <=  32'b00111111010010110001000101101101 ;
        2689:  q   <=  32'b00111111011101011001110111010100 ;
        2690:  q   <=  32'b00111111100010110010011000101111 ;
        2691:  q   <=  32'b00111111001001011010110011011001 ;
        2692:  q   <=  32'b00111111001000011110111011001110 ;
        2693:  q   <=  32'b00111111111100111001111010001110 ;
        2694:  q   <=  32'b10111111100101000111101110110111 ;
        2695:  q   <=  32'b10111110101100011101001010000101 ;
        2696:  q   <=  32'b10111111110110001111011111100000 ;
        2697:  q   <=  32'b00111111011010110101110011100010 ;
        2698:  q   <=  32'b00111100101100000110001000111100 ;
        2699:  q   <=  32'b10111110100110010100001100100010 ;
        2700:  q   <=  32'b10111111110111000100101000111111 ;
        2701:  q   <=  32'b00111110001110111101010110010000 ;
        2702:  q   <=  32'b10111110100001001111101110100001 ;
        2703:  q   <=  32'b10111111101011010110100110111001 ;
        2704:  q   <=  32'b10111111100101000010011100001111 ;
        2705:  q   <=  32'b10111111010000110001000110001001 ;
        2706:  q   <=  32'b10111110100000000010011101000100 ;
        2707:  q   <=  32'b10111111110100110000101010101011 ;
        2708:  q   <=  32'b10111110001110100101101110111111 ;
        2709:  q   <=  32'b00111111000111011001110110101101 ;
        2710:  q   <=  32'b10111110110000001101101101110011 ;
        2711:  q   <=  32'b10111111001100101011001001110000 ;
        2712:  q   <=  32'b00111110100110111011010111101111 ;
        2713:  q   <=  32'b00111111100011001111000000101111 ;
        2714:  q   <=  32'b10111110111001001010100111001100 ;
        2715:  q   <=  32'b10111110111011101111010011101000 ;
        2716:  q   <=  32'b10111111101101111100100011111000 ;
        2717:  q   <=  32'b10111111011110100100101110011010 ;
        2718:  q   <=  32'b00111111000110110001101111101000 ;
        2719:  q   <=  32'b10111101111010001100001110110100 ;
        2720:  q   <=  32'b00111111010000111011101001001110 ;
        2721:  q   <=  32'b00111111001010110111111001100110 ;
        2722:  q   <=  32'b00111110110000000110011010111000 ;
        2723:  q   <=  32'b00111111010001000100001101011011 ;
        2724:  q   <=  32'b00111111110000110000000100100000 ;
        2725:  q   <=  32'b00111111000100111010101011000000 ;
        2726:  q   <=  32'b00111110110110100001100100100010 ;
        2727:  q   <=  32'b10111101001011111101100001100010 ;
        2728:  q   <=  32'b10111111100111110000001001111001 ;
        2729:  q   <=  32'b10111111000000010100010010000011 ;
        2730:  q   <=  32'b00111110101001101101010111111011 ;
        2731:  q   <=  32'b10111111100011100100001100011110 ;
        2732:  q   <=  32'b00111110111011111011010111011011 ;
        2733:  q   <=  32'b00111110101001010010110110000011 ;
        2734:  q   <=  32'b00111101110011001101100000001010 ;
        2735:  q   <=  32'b00111110100110100101010110100010 ;
        2736:  q   <=  32'b00111100110000110010100111001010 ;
        2737:  q   <=  32'b10111100101101001010110000100001 ;
        2738:  q   <=  32'b10111100000011110111110101101010 ;
        2739:  q   <=  32'b00111111011011011111000011000101 ;
        2740:  q   <=  32'b10111101101110010011010010010011 ;
        2741:  q   <=  32'b11000000001010010000100010001000 ;
        2742:  q   <=  32'b10111110111110001110100010100110 ;
        2743:  q   <=  32'b00111110010010001010110001000010 ;
        2744:  q   <=  32'b00111111011101011011000001011010 ;
        2745:  q   <=  32'b00111111101100001010111001111000 ;
        2746:  q   <=  32'b10111111011100010000001111000010 ;
        2747:  q   <=  32'b00111111010000101100100001000000 ;
        2748:  q   <=  32'b00111110011100111010000101101010 ;
        2749:  q   <=  32'b10111110010101010101111111011010 ;
        2750:  q   <=  32'b00111100110010101010100111011100 ;
        2751:  q   <=  32'b10111100111001100001111101010000 ;
        2752:  q   <=  32'b00111110000011111011101001001101 ;
        2753:  q   <=  32'b00111110011100110100100111001010 ;
        2754:  q   <=  32'b10111111001010111110101010011110 ;
        2755:  q   <=  32'b10111111100001011100001010001111 ;
        2756:  q   <=  32'b00111111011101110011110001111011 ;
        2757:  q   <=  32'b10111110011000010000011111011010 ;
        2758:  q   <=  32'b00111111101101010000111110000010 ;
        2759:  q   <=  32'b10111111011011001001011101111111 ;
        2760:  q   <=  32'b10111111000110000001100110011100 ;
        2761:  q   <=  32'b00111111101101011110110001011010 ;
        2762:  q   <=  32'b00111111101101000010110001111100 ;
        2763:  q   <=  32'b10111111100000111011011001001011 ;
        2764:  q   <=  32'b00111110010100110111011111110001 ;
        2765:  q   <=  32'b00111111101010111010100110001001 ;
        2766:  q   <=  32'b00111111101010101001011001110100 ;
        2767:  q   <=  32'b10111111101001000111011101101101 ;
        2768:  q   <=  32'b00111111110011110010011011110000 ;
        2769:  q   <=  32'b00111111001010010110000101111100 ;
        2770:  q   <=  32'b00111110011010001100110110000001 ;
        2771:  q   <=  32'b10111110011001101111110101101101 ;
        2772:  q   <=  32'b10111111011101110100101101011000 ;
        2773:  q   <=  32'b00111101110000101001100010111001 ;
        2774:  q   <=  32'b10111110100000110111001001110001 ;
        2775:  q   <=  32'b01000000000100111101100100110001 ;
        2776:  q   <=  32'b00111110010000101001111100000100 ;
        2777:  q   <=  32'b10111110001100011001000011010001 ;
        2778:  q   <=  32'b10111100011001011101100100100110 ;
        2779:  q   <=  32'b10111111000111001101110001101011 ;
        2780:  q   <=  32'b01000000000001001001100001011110 ;
        2781:  q   <=  32'b00111111001000110001010000000010 ;
        2782:  q   <=  32'b00111101100110010110000111111101 ;
        2783:  q   <=  32'b00111111100011111100011100111000 ;
        2784:  q   <=  32'b10111101000001111011000100101001 ;
        2785:  q   <=  32'b10111101110010000010111111110010 ;
        2786:  q   <=  32'b10111111000011100111111010100100 ;
        2787:  q   <=  32'b10111111000111011001000101010111 ;
        2788:  q   <=  32'b00111111110011010110000111111111 ;
        2789:  q   <=  32'b00111111010001001011110000011101 ;
        2790:  q   <=  32'b00111101101100100000101000101101 ;
        2791:  q   <=  32'b00111111110110100010100001110000 ;
        2792:  q   <=  32'b00111100110000011001101111001001 ;
        2793:  q   <=  32'b00111110100101001000000001111110 ;
        2794:  q   <=  32'b10111111101101011011111101000001 ;
        2795:  q   <=  32'b00111110111100110101011100001110 ;
        2796:  q   <=  32'b10111111101110010100000111000000 ;
        2797:  q   <=  32'b10111111011111001111111111101010 ;
        2798:  q   <=  32'b00111111011100110000101010001001 ;
        2799:  q   <=  32'b00111110101100111101001110100000 ;
        2800:  q   <=  32'b10111111010111110100110111011000 ;
        2801:  q   <=  32'b10111110110010111101011101010011 ;
        2802:  q   <=  32'b00111110100000110100101110010000 ;
        2803:  q   <=  32'b00111110011000010100111001011010 ;
        2804:  q   <=  32'b10111111110110110001000001111100 ;
        2805:  q   <=  32'b10111111100110100101011000110000 ;
        2806:  q   <=  32'b10111111111000101110111011010101 ;
        2807:  q   <=  32'b10111101100101000111011001111111 ;
        2808:  q   <=  32'b10111111110111000100110101111101 ;
        2809:  q   <=  32'b00111111001100111010111001111100 ;
        2810:  q   <=  32'b10111111100000001011001100101100 ;
        2811:  q   <=  32'b10111111100011011001111101100100 ;
        2812:  q   <=  32'b00111111111001010011000100010001 ;
        2813:  q   <=  32'b01000000000010100110010010000000 ;
        2814:  q   <=  32'b10111111010100011011110000101011 ;
        2815:  q   <=  32'b10111101000101111100000101001111 ;
        2816:  q   <=  32'b00111111111110110100001110110110 ;
        2817:  q   <=  32'b10111111000010100100111011100101 ;
        2818:  q   <=  32'b00111111110110111101011100101010 ;
        2819:  q   <=  32'b00111111010100011101111011110100 ;
        2820:  q   <=  32'b00111101011000110110100111010000 ;
        2821:  q   <=  32'b10111110101101001100110011011000 ;
        2822:  q   <=  32'b00111111110110001011100100011101 ;
        2823:  q   <=  32'b00111111001101100000011101100110 ;
        2824:  q   <=  32'b10111111001000011111110011010001 ;
        2825:  q   <=  32'b00111110110010010001001101101110 ;
        2826:  q   <=  32'b10111111011000001100001000010110 ;
        2827:  q   <=  32'b00111110000110001000010100100110 ;
        2828:  q   <=  32'b00111111110001000001010010010100 ;
        2829:  q   <=  32'b00111111000010000010011100101100 ;
        2830:  q   <=  32'b10111111010000100111100110001011 ;
        2831:  q   <=  32'b00111110101100100010101011111010 ;
        2832:  q   <=  32'b10111111001100101010001100110010 ;
        2833:  q   <=  32'b01000000000000010011110001110100 ;
        2834:  q   <=  32'b10111111111001011001011111110010 ;
        2835:  q   <=  32'b10111111001010001101010101111100 ;
        2836:  q   <=  32'b00111111010001010111110111110111 ;
        2837:  q   <=  32'b10111111010100100000000111011111 ;
        2838:  q   <=  32'b00111100100100101000101000111100 ;
        2839:  q   <=  32'b00111111001001111000111110011110 ;
        2840:  q   <=  32'b00111111101000001111110001000101 ;
        2841:  q   <=  32'b10111111011011010101010100011101 ;
        2842:  q   <=  32'b10111110001011011111010001101001 ;
        2843:  q   <=  32'b10111110111100010111111100001110 ;
        2844:  q   <=  32'b10111101111010011111001100111111 ;
        2845:  q   <=  32'b00111110101111010010110101100010 ;
        2846:  q   <=  32'b10111111000111100101110110010010 ;
        2847:  q   <=  32'b00111111010011001101010001011000 ;
        2848:  q   <=  32'b00111110110110100111011111100111 ;
        2849:  q   <=  32'b10111110111100011101010101010110 ;
        2850:  q   <=  32'b00111110100011010100100110001101 ;
        2851:  q   <=  32'b00111111011110111111011001001110 ;
        2852:  q   <=  32'b00111111011111100011110001001001 ;
        2853:  q   <=  32'b00111111001010110000111111000000 ;
        2854:  q   <=  32'b10111101100001010001110111100100 ;
        2855:  q   <=  32'b10111111000111101011111011001000 ;
        2856:  q   <=  32'b00111110011001010111101110010110 ;
        2857:  q   <=  32'b10111110111011101010100101100111 ;
        2858:  q   <=  32'b10111110101010100000011101001010 ;
        2859:  q   <=  32'b00111111011011001100000010101001 ;
        2860:  q   <=  32'b00111111101110010011100000100001 ;
        2861:  q   <=  32'b00111111000110001000100001110011 ;
        2862:  q   <=  32'b01000000000000110110100011001000 ;
        2863:  q   <=  32'b10111111110000111011111001111001 ;
        2864:  q   <=  32'b00111100101110011101101101001011 ;
        2865:  q   <=  32'b00111101110000110010010010101110 ;
        2866:  q   <=  32'b00111111110011101010100011001100 ;
        2867:  q   <=  32'b00111111000000000101001101110000 ;
        2868:  q   <=  32'b10111110101001011100111001100010 ;
        2869:  q   <=  32'b00111111000011011110000100100011 ;
        2870:  q   <=  32'b00111111001001000111011100101100 ;
        2871:  q   <=  32'b00111110001110110000001000010011 ;
        2872:  q   <=  32'b11000000000000011100001000101100 ;
        2873:  q   <=  32'b00111111100000101111010001010000 ;
        2874:  q   <=  32'b11000000010111110111010101101011 ;
        2875:  q   <=  32'b00111101111000000011110000011010 ;
        2876:  q   <=  32'b10111111110001101001001000000111 ;
        2877:  q   <=  32'b10111110101101011101000100011000 ;
        2878:  q   <=  32'b00111111101100110000001111101110 ;
        2879:  q   <=  32'b10111111000000110111001100011000 ;
        2880:  q   <=  32'b00111111111101010110011000100100 ;
        2881:  q   <=  32'b00111111010001110100010111101010 ;
        2882:  q   <=  32'b10111110011111000101111010111010 ;
        2883:  q   <=  32'b10111111011001110100110111011001 ;
        2884:  q   <=  32'b10111110111111011110011011100110 ;
        2885:  q   <=  32'b00111110101111111011110111000111 ;
        2886:  q   <=  32'b11000000000101111011011011001100 ;
        2887:  q   <=  32'b00111111000111010111010010110100 ;
        2888:  q   <=  32'b00111110100011110001011000001000 ;
        2889:  q   <=  32'b00111111010100011010000100100100 ;
        2890:  q   <=  32'b01000000000000110000101001011000 ;
        2891:  q   <=  32'b10111110101001011100000111010001 ;
        2892:  q   <=  32'b10111111011110110000010011010001 ;
        2893:  q   <=  32'b00111111100101101111111001000000 ;
        2894:  q   <=  32'b00111111011001010000001101100000 ;
        2895:  q   <=  32'b10111110000100100101110001100111 ;
        2896:  q   <=  32'b10111111000101111110110110101111 ;
        2897:  q   <=  32'b00111110011111101110010000100110 ;
        2898:  q   <=  32'b10111111100100001001110010110101 ;
        2899:  q   <=  32'b00111101100001110101110010011100 ;
        2900:  q   <=  32'b10111111001000110100111100000110 ;
        2901:  q   <=  32'b10111111010100011011111000100101 ;
        2902:  q   <=  32'b00111111011101111100101111001101 ;
        2903:  q   <=  32'b00111100111110001001111001111100 ;
        2904:  q   <=  32'b00111111101011001111000010111011 ;
        2905:  q   <=  32'b10111111100010110000111001001111 ;
        2906:  q   <=  32'b00111110011101100000100000001001 ;
        2907:  q   <=  32'b10111111100001011110100101000100 ;
        2908:  q   <=  32'b00111111000111100110010001000111 ;
        2909:  q   <=  32'b00111111101001110000101101011100 ;
        2910:  q   <=  32'b00111111100000110000000111000001 ;
        2911:  q   <=  32'b11000000000001110110001001101101 ;
        2912:  q   <=  32'b00111111001011101000010111001000 ;
        2913:  q   <=  32'b00111100000011101011000101011001 ;
        2914:  q   <=  32'b00111110101010110010010111011111 ;
        2915:  q   <=  32'b10111111000011000010001100111110 ;
        2916:  q   <=  32'b10111111110100110101001101110100 ;
        2917:  q   <=  32'b00111111011001001000111000011001 ;
        2918:  q   <=  32'b10111111000000011100111001100100 ;
        2919:  q   <=  32'b10111110101010001101101001100010 ;
        2920:  q   <=  32'b00111110001011000110010011110000 ;
        2921:  q   <=  32'b01000000001000100101100111110010 ;
        2922:  q   <=  32'b01000000000100101100101011000111 ;
        2923:  q   <=  32'b10111111101010001100100111100001 ;
        2924:  q   <=  32'b10111110111100101100000111001001 ;
        2925:  q   <=  32'b00111111011111001100010100010000 ;
        2926:  q   <=  32'b11000000000001001010110001110111 ;
        2927:  q   <=  32'b00111111100111110011110000111111 ;
        2928:  q   <=  32'b10111110101000010110011100010101 ;
        2929:  q   <=  32'b00111111101100110001110000010000 ;
        2930:  q   <=  32'b10111111011000010011111111101000 ;
        2931:  q   <=  32'b10111111011011000010011100100111 ;
        2932:  q   <=  32'b01000000000101000001111100101101 ;
        2933:  q   <=  32'b00111111000101101000100000001000 ;
        2934:  q   <=  32'b10111110100111101001100111011101 ;
        2935:  q   <=  32'b10111111100001000011100000101011 ;
        2936:  q   <=  32'b00111111100011010011101010011000 ;
        2937:  q   <=  32'b00111110101011110010100011100110 ;
        2938:  q   <=  32'b11000000000100001110010101000011 ;
        2939:  q   <=  32'b10111111011001110011110110111101 ;
        2940:  q   <=  32'b01000000001111100001010011110100 ;
        2941:  q   <=  32'b10111100010000001100011101101100 ;
        2942:  q   <=  32'b10111111111111111111000011100101 ;
        2943:  q   <=  32'b10111111011000110101010011111000 ;
        2944:  q   <=  32'b10111110110101101111110101110010 ;
        2945:  q   <=  32'b00111111001100011100111111100011 ;
        2946:  q   <=  32'b10111110001001101010100010100100 ;
        2947:  q   <=  32'b00111101110100000000011101101010 ;
        2948:  q   <=  32'b10111100100100100100101111101000 ;
        2949:  q   <=  32'b10111111011101011101011111111111 ;
        2950:  q   <=  32'b00111111100101100001111001111110 ;
        2951:  q   <=  32'b10111110101110110000010100000101 ;
        2952:  q   <=  32'b10111110111011010100010000101000 ;
        2953:  q   <=  32'b00111110010001111010101101011000 ;
        2954:  q   <=  32'b10111101100010010001101100111111 ;
        2955:  q   <=  32'b10111111000001011000001011111111 ;
        2956:  q   <=  32'b00111110000000100010011001110000 ;
        2957:  q   <=  32'b01000000000001110011101110110001 ;
        2958:  q   <=  32'b00111111000010101001000101100101 ;
        2959:  q   <=  32'b10111111001001111011001110101011 ;
        2960:  q   <=  32'b10111111010111101001100101101111 ;
        2961:  q   <=  32'b10111110011101001010000110100110 ;
        2962:  q   <=  32'b10111111110010011011100111110011 ;
        2963:  q   <=  32'b00111111111010011011001000110111 ;
        2964:  q   <=  32'b00111110010100010010101101111110 ;
        2965:  q   <=  32'b10111111100101001110101000100111 ;
        2966:  q   <=  32'b00111101111101110000001001000111 ;
        2967:  q   <=  32'b10111111101110001100010100110101 ;
        2968:  q   <=  32'b00111111000101010001010010100001 ;
        2969:  q   <=  32'b10111110001110011101001000010101 ;
        2970:  q   <=  32'b00111101001011000001001001110010 ;
        2971:  q   <=  32'b00111110101110010100001101011000 ;
        2972:  q   <=  32'b00111111010110101000110100001010 ;
        2973:  q   <=  32'b10111111010011110100110100111000 ;
        2974:  q   <=  32'b10111111101110111100100001010000 ;
        2975:  q   <=  32'b10111101110101001100011110001100 ;
        2976:  q   <=  32'b10111111010100101010101001110011 ;
        2977:  q   <=  32'b00111110110110011001011100101010 ;
        2978:  q   <=  32'b10111111111011010110011001001100 ;
        2979:  q   <=  32'b00111111010110111100101110010011 ;
        2980:  q   <=  32'b00111110100111001101111110100000 ;
        2981:  q   <=  32'b10111111100011100100011110100111 ;
        2982:  q   <=  32'b10111110101000100110110101100000 ;
        2983:  q   <=  32'b00111111010101100111111000101010 ;
        2984:  q   <=  32'b01000000000110110100101100110101 ;
        2985:  q   <=  32'b10111110101100111100000111111110 ;
        2986:  q   <=  32'b00111111101100001110010000100000 ;
        2987:  q   <=  32'b10111111010111000101001111101010 ;
        2988:  q   <=  32'b00111110010100111101101100011000 ;
        2989:  q   <=  32'b10111110010101000111101000100111 ;
        2990:  q   <=  32'b00111110101011100011011000101011 ;
        2991:  q   <=  32'b10111110111111110000100010001110 ;
        2992:  q   <=  32'b10111111101101011111000001000010 ;
        2993:  q   <=  32'b10111110100010101010001011101000 ;
        2994:  q   <=  32'b00111110111000010001101110000101 ;
        2995:  q   <=  32'b10111111000000011001001010100011 ;
        2996:  q   <=  32'b10111110001111001100010111001000 ;
        2997:  q   <=  32'b00111110110011011101001011010000 ;
        2998:  q   <=  32'b00111111000010100000101011011100 ;
        2999:  q   <=  32'b10111111001110111100110011000011 ;
        3000:  q   <=  32'b10111110100010010110100000001101 ;
        3001:  q   <=  32'b00111111010111101101111110001001 ;
        3002:  q   <=  32'b00111110101010010101100101110001 ;
        3003:  q   <=  32'b10111111101011001000011111100000 ;
        3004:  q   <=  32'b00111111110001100010000010101001 ;
        3005:  q   <=  32'b10111111000111011101101111100111 ;
        3006:  q   <=  32'b10111111001100101101010110001011 ;
        3007:  q   <=  32'b10111111101101100011100001011101 ;
        3008:  q   <=  32'b10111101111000001000011011101110 ;
        3009:  q   <=  32'b10111101110100100101101010111001 ;
        3010:  q   <=  32'b10111110101001010011101100011100 ;
        3011:  q   <=  32'b10111111010101101110111100110010 ;
        3012:  q   <=  32'b10111111110101001000110011101111 ;
        3013:  q   <=  32'b01000000010000001100110010010100 ;
        3014:  q   <=  32'b00111111110000000001101110001010 ;
        3015:  q   <=  32'b10111110101101111100110111000000 ;
        3016:  q   <=  32'b10111101111010110100010111011010 ;
        3017:  q   <=  32'b00111110101101111100000111100100 ;
        3018:  q   <=  32'b10111100010001101101101111000001 ;
        3019:  q   <=  32'b10111111000100100000001100011000 ;
        3020:  q   <=  32'b00111111011011110001110011100111 ;
        3021:  q   <=  32'b10111111100100011011010001011101 ;
        3022:  q   <=  32'b00111111111110101000011011000111 ;
        3023:  q   <=  32'b10111111111000011011000110000000 ;
        3024:  q   <=  32'b10111110101001011000110000010011 ;
        3025:  q   <=  32'b00111111010111110110001000110011 ;
        3026:  q   <=  32'b00111101111100010111110110011111 ;
        3027:  q   <=  32'b10111111110000000110010000011001 ;
        3028:  q   <=  32'b00111111011010111111110101100100 ;
        3029:  q   <=  32'b00111110001001110010100110101100 ;
        3030:  q   <=  32'b10111111010100001000111001000100 ;
        3031:  q   <=  32'b00111110110011101011001100010110 ;
        3032:  q   <=  32'b00111111010000011001001110001000 ;
        3033:  q   <=  32'b01000000000010111100110111011100 ;
        3034:  q   <=  32'b10111101110000000001000100001111 ;
        3035:  q   <=  32'b10111110100101101010001000101110 ;
        3036:  q   <=  32'b10111111000000010011101011110000 ;
        3037:  q   <=  32'b10111111111101101010011111100111 ;
        3038:  q   <=  32'b00111111000001010111100100110100 ;
        3039:  q   <=  32'b11000000000000110111101101111001 ;
        3040:  q   <=  32'b10111110100010100010100000100100 ;
        3041:  q   <=  32'b10111110100011001101000100000000 ;
        3042:  q   <=  32'b00111111010110000101101101101000 ;
        3043:  q   <=  32'b11000000001100010101101100001001 ;
        3044:  q   <=  32'b00111111011010110000011011110101 ;
        3045:  q   <=  32'b10111111000001001110110111011010 ;
        3046:  q   <=  32'b10111111101001011000000101101100 ;
        3047:  q   <=  32'b10111100000011101101011001010100 ;
        3048:  q   <=  32'b00111110011011101111010000000001 ;
        3049:  q   <=  32'b10111110110110010011000000101101 ;
        3050:  q   <=  32'b10111111101111000001011011100100 ;
        3051:  q   <=  32'b00111111100110100110101111111011 ;
        3052:  q   <=  32'b00111110010010100001010000010100 ;
        3053:  q   <=  32'b10111111001101001111010111001011 ;
        3054:  q   <=  32'b00111111100110111011000111101100 ;
        3055:  q   <=  32'b00111110101110111111110111000010 ;
        3056:  q   <=  32'b10111111101000100011110111110011 ;
        3057:  q   <=  32'b00111111000111101111110100100011 ;
        3058:  q   <=  32'b10111111111001011101000101110100 ;
        3059:  q   <=  32'b10111111100001110110011101001000 ;
        3060:  q   <=  32'b00111110000110110010111001111001 ;
        3061:  q   <=  32'b00111110110100101001000100110100 ;
        3062:  q   <=  32'b00111101100100000110000100100100 ;
        3063:  q   <=  32'b10111111111101110110110101101010 ;
        3064:  q   <=  32'b00111111010100011001011111000100 ;
        3065:  q   <=  32'b00111111101000011000000101000001 ;
        3066:  q   <=  32'b00111111100101010110101101111101 ;
        3067:  q   <=  32'b10111111000100100000000100100101 ;
        3068:  q   <=  32'b10111110110010011010110011110001 ;
        3069:  q   <=  32'b10111111100000100011101101000111 ;
        3070:  q   <=  32'b00111110100000000001101011111011 ;
        3071:  q   <=  32'b00111110100000010001011010000000 ;
        3072:  q   <=  32'b10111111010001010111111110100100 ;
        3073:  q   <=  32'b00111111011010110110011101010100 ;
        3074:  q   <=  32'b00111111010110100010011011111111 ;
        3075:  q   <=  32'b00111111001010000011100101101100 ;
        3076:  q   <=  32'b10111111010000001110001100001001 ;
        3077:  q   <=  32'b10111111101010110101010000000111 ;
        3078:  q   <=  32'b00111111001001101111100000111001 ;
        3079:  q   <=  32'b00111111101110010011111001100101 ;
        3080:  q   <=  32'b10111111101001010010001011011001 ;
        3081:  q   <=  32'b11000000000011010101001011111000 ;
        3082:  q   <=  32'b00111111101101111101001001100100 ;
        3083:  q   <=  32'b10111101011111001001101111111101 ;
        3084:  q   <=  32'b00111111100101101100001001011100 ;
        3085:  q   <=  32'b00111111011111000100101010011011 ;
        3086:  q   <=  32'b10111111100110111111101001100000 ;
        3087:  q   <=  32'b10111110110111010001111100100110 ;
        3088:  q   <=  32'b10111111010101011011111010110110 ;
        3089:  q   <=  32'b00111110001101111111111000001111 ;
        3090:  q   <=  32'b00111111100101010100100101100101 ;
        3091:  q   <=  32'b00111101011001010101000110000011 ;
        3092:  q   <=  32'b11000000000001100110011100010101 ;
        3093:  q   <=  32'b00111111100111100001111000110111 ;
        3094:  q   <=  32'b00111011001011110001010011001001 ;
        3095:  q   <=  32'b10111110111010110100100001101000 ;
        3096:  q   <=  32'b11000000000001101001101001110001 ;
        3097:  q   <=  32'b00111110101111110111001010101001 ;
        3098:  q   <=  32'b00111110011110110001000010011001 ;
        3099:  q   <=  32'b00111110101011010101101001000000 ;
        3100:  q   <=  32'b10111111100010011111111000001010 ;
        3101:  q   <=  32'b10111111001110101110101111101011 ;
        3102:  q   <=  32'b10111111011010101001010001101100 ;
        3103:  q   <=  32'b00111111111001001100111010001010 ;
        3104:  q   <=  32'b10111111010100100000010111110111 ;
        3105:  q   <=  32'b10111110010010010110111010110010 ;
        3106:  q   <=  32'b10111111011000111110000001110101 ;
        3107:  q   <=  32'b00111111011010010010011011010010 ;
        3108:  q   <=  32'b10111100010010001111010000101111 ;
        3109:  q   <=  32'b00111101100101010001111111000010 ;
        3110:  q   <=  32'b00111111011100000111110110010110 ;
        3111:  q   <=  32'b00111111001011001101110001011010 ;
        3112:  q   <=  32'b00111111010010010011010100111011 ;
        3113:  q   <=  32'b11000000000010000111111011010010 ;
        3114:  q   <=  32'b00111110011000010011010100111100 ;
        3115:  q   <=  32'b00111111011101110101111001111101 ;
        3116:  q   <=  32'b00111110101100110011001001101101 ;
        3117:  q   <=  32'b00111111011001101101110101011101 ;
        3118:  q   <=  32'b01000000000001111100000110001101 ;
        3119:  q   <=  32'b00111111100111111101000110110000 ;
        3120:  q   <=  32'b10111111100011111100010010001101 ;
        3121:  q   <=  32'b10111111010101001000000001110100 ;
        3122:  q   <=  32'b10111101111110010110011100100001 ;
        3123:  q   <=  32'b10111111001001001000000011011000 ;
        3124:  q   <=  32'b10111101101000011011000010000101 ;
        3125:  q   <=  32'b00111111100111010011001011001100 ;
        3126:  q   <=  32'b10111111000010000000011110010111 ;
        3127:  q   <=  32'b10111110100100100111110001010100 ;
        3128:  q   <=  32'b10111110011010010001000101110100 ;
        3129:  q   <=  32'b00111111001011001010110110001100 ;
        3130:  q   <=  32'b00111111100001001011011100101100 ;
        3131:  q   <=  32'b10111110000110010000110010110100 ;
        3132:  q   <=  32'b10111110101000100101100001111100 ;
        3133:  q   <=  32'b00111111011011110000000000001111 ;
        3134:  q   <=  32'b00111111001110010010100100100101 ;
        3135:  q   <=  32'b00111110111110011111001101011100 ;
        3136:  q   <=  32'b01000000010100010000100101100110 ;
        3137:  q   <=  32'b00111101000000011101100010100111 ;
        3138:  q   <=  32'b00111110101011101011101110010110 ;
        3139:  q   <=  32'b10111101101010110001001001001011 ;
        3140:  q   <=  32'b00111111000111011100110111000101 ;
        3141:  q   <=  32'b10111111000001100110011001011000 ;
        3142:  q   <=  32'b00111111100000001111110010001000 ;
        3143:  q   <=  32'b00111111111010100010000000000101 ;
        3144:  q   <=  32'b00111101101011101010101110000010 ;
        3145:  q   <=  32'b10111101100010111110110111010101 ;
        3146:  q   <=  32'b10111111000100000011111101000100 ;
        3147:  q   <=  32'b10111110111100100111100001001100 ;
        3148:  q   <=  32'b10111111110110100000110101101011 ;
        3149:  q   <=  32'b10111101010111000000100110001101 ;
        3150:  q   <=  32'b10111111011000011001111111000011 ;
        3151:  q   <=  32'b00111111101000001100000100001100 ;
        3152:  q   <=  32'b00111110000111111001010011101101 ;
        3153:  q   <=  32'b00111101011000010000000100010111 ;
        3154:  q   <=  32'b00111111101100110000001111000100 ;
        3155:  q   <=  32'b10111111111000110100100001110010 ;
        3156:  q   <=  32'b00111110101010001100100001101010 ;
        3157:  q   <=  32'b10111111100001110110100101011011 ;
        3158:  q   <=  32'b10111111001001001011001111010111 ;
        3159:  q   <=  32'b00111110100001000101001001011001 ;
        3160:  q   <=  32'b00111111011001000100011000010011 ;
        3161:  q   <=  32'b10111111010101100010110011100010 ;
        3162:  q   <=  32'b00111111000011011001101100011111 ;
        3163:  q   <=  32'b00111111101110101010110100101000 ;
        3164:  q   <=  32'b10111111010110101110011010101010 ;
        3165:  q   <=  32'b10111111011111011111101110111111 ;
        3166:  q   <=  32'b10111100001111111010111011101001 ;
        3167:  q   <=  32'b00111111001000000111110100111000 ;
        3168:  q   <=  32'b00111010110001001000000101100000 ;
        3169:  q   <=  32'b10111111010100001111101011001010 ;
        3170:  q   <=  32'b00111101111010111101001001111000 ;
        3171:  q   <=  32'b00111110010101000000100111001110 ;
        3172:  q   <=  32'b10111110111000111001110110011010 ;
        3173:  q   <=  32'b10111111100011110110110000110101 ;
        3174:  q   <=  32'b00111110110111101110011100111101 ;
        3175:  q   <=  32'b00111100100010111111110101110110 ;
        3176:  q   <=  32'b10111110101110011101100101000000 ;
        3177:  q   <=  32'b10111111001000011001100011000111 ;
        3178:  q   <=  32'b10111111000000000001010101001100 ;
        3179:  q   <=  32'b10111111010111100000000001011111 ;
        3180:  q   <=  32'b10111111100001010010000111000101 ;
        3181:  q   <=  32'b00111111101000011111100110101000 ;
        3182:  q   <=  32'b10111110011101110100000010111010 ;
        3183:  q   <=  32'b10111111110111010101000011100110 ;
        3184:  q   <=  32'b10111110111110011111101010110101 ;
        3185:  q   <=  32'b00111111100001111011101010101100 ;
        3186:  q   <=  32'b10111111000010011100010001110101 ;
        3187:  q   <=  32'b00111111111000110111111111001101 ;
        3188:  q   <=  32'b10111111010001111000111010001011 ;
        3189:  q   <=  32'b10111111010000001100001011000100 ;
        3190:  q   <=  32'b10111111100001000011110110110110 ;
        3191:  q   <=  32'b00111111100101001111100010101001 ;
        3192:  q   <=  32'b10111111000101001000000111010100 ;
        3193:  q   <=  32'b00111110110101011010100010101000 ;
        3194:  q   <=  32'b10111111110100101111010111000010 ;
        3195:  q   <=  32'b10111111000100101001101011011011 ;
        3196:  q   <=  32'b00111111001010001100001101101110 ;
        3197:  q   <=  32'b10111111101000111110010000110011 ;
        3198:  q   <=  32'b00111101010011010100111011100000 ;
        3199:  q   <=  32'b00111111000011000110010000100010 ;
        3200:  q   <=  32'b00111111111000111010010000100100 ;
        3201:  q   <=  32'b00111111001001000001111001001010 ;
        3202:  q   <=  32'b00111111011100100101101100100111 ;
        3203:  q   <=  32'b10111110101101010110000011101001 ;
        3204:  q   <=  32'b10111111000101000010110101011100 ;
        3205:  q   <=  32'b00111101011001110101000010010000 ;
        3206:  q   <=  32'b10111111011001001011000011001011 ;
        3207:  q   <=  32'b00111111100011111010000000111111 ;
        3208:  q   <=  32'b00111111010001101001110010110110 ;
        3209:  q   <=  32'b00111111011101100110011000011100 ;
        3210:  q   <=  32'b00111111101000010110000101011111 ;
        3211:  q   <=  32'b10111101110111010000010001100010 ;
        3212:  q   <=  32'b10111111000100111100000010011000 ;
        3213:  q   <=  32'b00111111000001101000111111011011 ;
        3214:  q   <=  32'b00111111100100110111001101101010 ;
        3215:  q   <=  32'b00111111010110111011111010110111 ;
        3216:  q   <=  32'b00111111011100100001000101001000 ;
        3217:  q   <=  32'b00111111110000001100100011100001 ;
        3218:  q   <=  32'b00111110100101110011011010001000 ;
        3219:  q   <=  32'b00111111100110100001111111011001 ;
        3220:  q   <=  32'b10111100010000100001010011101001 ;
        3221:  q   <=  32'b00111111010010100001110010110001 ;
        3222:  q   <=  32'b10111111101100111010100010010100 ;
        3223:  q   <=  32'b00111111110001010110001110111011 ;
        3224:  q   <=  32'b10111111111000110011000000100101 ;
        3225:  q   <=  32'b00111110010100101001011110100000 ;
        3226:  q   <=  32'b10111110101100010100001001101100 ;
        3227:  q   <=  32'b10111111100101000101100110001100 ;
        3228:  q   <=  32'b00111110101010111111000101101101 ;
        3229:  q   <=  32'b00111110101010100001101111000011 ;
        3230:  q   <=  32'b00111111101101001010001010000010 ;
        3231:  q   <=  32'b00111110000011000010010111001011 ;
        3232:  q   <=  32'b00111111000100111101111101101111 ;
        3233:  q   <=  32'b00111110011110001110110000001110 ;
        3234:  q   <=  32'b00111111101110111101110010100101 ;
        3235:  q   <=  32'b00111111100100001011010111111110 ;
        3236:  q   <=  32'b00111100001011101000101010011000 ;
        3237:  q   <=  32'b00111101111111101010001010101001 ;
        3238:  q   <=  32'b00111111111000111100010001100110 ;
        3239:  q   <=  32'b10111110011101010011100000110111 ;
        3240:  q   <=  32'b00111111010110111010010101100101 ;
        3241:  q   <=  32'b10111111011000001101101111011011 ;
        3242:  q   <=  32'b10111111010000110000111011100100 ;
        3243:  q   <=  32'b00111111010111001101111101010011 ;
        3244:  q   <=  32'b00111111001001011111011101010011 ;
        3245:  q   <=  32'b00111111100001110110111110010001 ;
        3246:  q   <=  32'b10111111001000100001100011010100 ;
        3247:  q   <=  32'b00111111100000100100110101111010 ;
        3248:  q   <=  32'b00111110001100000000110101001000 ;
        3249:  q   <=  32'b10111101010000100111010000110000 ;
        3250:  q   <=  32'b00111111110110000011010111101011 ;
        3251:  q   <=  32'b00111111101101111111000100010010 ;
        3252:  q   <=  32'b11000000000100000001000110101010 ;
        3253:  q   <=  32'b00111110101101101000010110111110 ;
        3254:  q   <=  32'b10111111010110011010100101101110 ;
        3255:  q   <=  32'b10111110100110010101111011000000 ;
        3256:  q   <=  32'b10111111001000100101111000011101 ;
        3257:  q   <=  32'b00111111110011111110111011011111 ;
        3258:  q   <=  32'b00111111100111101101101101100010 ;
        3259:  q   <=  32'b00111111000011100010011011011101 ;
        3260:  q   <=  32'b00111111001101000001001100101101 ;
        3261:  q   <=  32'b00111110111010101001010001100010 ;
        3262:  q   <=  32'b00111111001011110001100110010011 ;
        3263:  q   <=  32'b00111110100000001010100100000111 ;
        3264:  q   <=  32'b10111110001101101100100110111001 ;
        3265:  q   <=  32'b00111111000000011111101001010001 ;
        3266:  q   <=  32'b10111110100111101010101100011000 ;
        3267:  q   <=  32'b10111110110010011110101011100101 ;
        3268:  q   <=  32'b10111110100010100001101100101011 ;
        3269:  q   <=  32'b10111101101101000111110110010111 ;
        3270:  q   <=  32'b00111100000000111000110100110111 ;
        3271:  q   <=  32'b01000000001000100000100011110000 ;
        3272:  q   <=  32'b10111111100111001001001100111010 ;
        3273:  q   <=  32'b10111111100010010010111100011111 ;
        3274:  q   <=  32'b00111110011110111111011011001100 ;
        3275:  q   <=  32'b10111101010011110100110111111010 ;
        3276:  q   <=  32'b10111111001110101110101100100110 ;
        3277:  q   <=  32'b00111110101001110110101011011011 ;
        3278:  q   <=  32'b00111111010000001100010000000011 ;
        3279:  q   <=  32'b10111111100100111010110100100101 ;
        3280:  q   <=  32'b10111110110100001101001111110011 ;
        3281:  q   <=  32'b10111111101001001101101000011110 ;
        3282:  q   <=  32'b00111101101010110010101011000111 ;
        3283:  q   <=  32'b00111110001001111011101100000000 ;
        3284:  q   <=  32'b00111111001011101011110100110111 ;
        3285:  q   <=  32'b10111111100010110000111000011000 ;
        3286:  q   <=  32'b00111110100110000101000011101011 ;
        3287:  q   <=  32'b10111110000100101011111101100110 ;
        3288:  q   <=  32'b00111111101100100010101110001001 ;
        3289:  q   <=  32'b00111110100111010000110111111101 ;
        3290:  q   <=  32'b10111111000010011000010011100111 ;
        3291:  q   <=  32'b10111110011010100110110100110110 ;
        3292:  q   <=  32'b10111111000010010100010110111101 ;
        3293:  q   <=  32'b00111111101110000011000111011001 ;
        3294:  q   <=  32'b10111111000000101101011101101101 ;
        3295:  q   <=  32'b10111111110011011010110011001000 ;
        3296:  q   <=  32'b10111110010011100001001010100110 ;
        3297:  q   <=  32'b00111111100100100101111001010001 ;
        3298:  q   <=  32'b00111111001010011100110101110001 ;
        3299:  q   <=  32'b00111110001010000000010110111011 ;
        3300:  q   <=  32'b00111111111001001000100000101010 ;
        3301:  q   <=  32'b10111111000101100111010001000010 ;
        3302:  q   <=  32'b00111110100001001010000001101000 ;
        3303:  q   <=  32'b10111111010111110011000001111011 ;
        3304:  q   <=  32'b10111111010010011011010011100101 ;
        3305:  q   <=  32'b10111110101100000100110101001100 ;
        3306:  q   <=  32'b00111111001001011100101000111011 ;
        3307:  q   <=  32'b01000000000000110111011011010000 ;
        3308:  q   <=  32'b00111111010011001000011101110010 ;
        3309:  q   <=  32'b10111111100010010001100100010000 ;
        3310:  q   <=  32'b10111110010100100001010001000111 ;
        3311:  q   <=  32'b10111111000011011110111111111011 ;
        3312:  q   <=  32'b10111110100101011111110010100011 ;
        3313:  q   <=  32'b00111111100101110001000111010111 ;
        3314:  q   <=  32'b00111110110000010011100111101101 ;
        3315:  q   <=  32'b00111111011111011101011111010001 ;
        3316:  q   <=  32'b00111111000110100111101111010010 ;
        3317:  q   <=  32'b10111111010010101111101010010101 ;
        3318:  q   <=  32'b00111111011011100100101000010111 ;
        3319:  q   <=  32'b10111111101011001101100110000110 ;
        3320:  q   <=  32'b00111111010011001011111100000000 ;
        3321:  q   <=  32'b00111111000110011000000111010110 ;
        3322:  q   <=  32'b00111111100011001101101011011010 ;
        3323:  q   <=  32'b10111111101101011011101000011001 ;
        3324:  q   <=  32'b10111110010100001000010111111010 ;
        3325:  q   <=  32'b00111100100100101011111001101100 ;
        3326:  q   <=  32'b00111101110011011000010100001110 ;
        3327:  q   <=  32'b00111111011000000101100011101000 ;
        3328:  q   <=  32'b00111111001100110110000010110010 ;
        3329:  q   <=  32'b00111111001001101110101010000001 ;
        3330:  q   <=  32'b00111110001101101101000010101011 ;
        3331:  q   <=  32'b00111111110101101000011110000010 ;
        3332:  q   <=  32'b10111110101001100111001100101011 ;
        3333:  q   <=  32'b00111101110011110010011010011000 ;
        3334:  q   <=  32'b10111111000100111010001000011010 ;
        3335:  q   <=  32'b10111101011111000000010011100110 ;
        3336:  q   <=  32'b00111111001110011100000000011110 ;
        3337:  q   <=  32'b10111111100111010001100110001001 ;
        3338:  q   <=  32'b00111110010000111000001101001111 ;
        3339:  q   <=  32'b10111111001111000001110100001110 ;
        3340:  q   <=  32'b00111111010010011101001110010001 ;
        3341:  q   <=  32'b10111111111110111001000110100101 ;
        3342:  q   <=  32'b10111111111110100100111010011110 ;
        3343:  q   <=  32'b00111111110011111110100011011001 ;
        3344:  q   <=  32'b10111110000110010000000110010010 ;
        3345:  q   <=  32'b10111111111110111111000000110101 ;
        3346:  q   <=  32'b10111111110101111101001101011010 ;
        3347:  q   <=  32'b10111101101100100000001111111111 ;
        3348:  q   <=  32'b00111110100111010110000110110101 ;
        3349:  q   <=  32'b00111110101011001101001011000111 ;
        3350:  q   <=  32'b00111111100010001001001100101111 ;
        3351:  q   <=  32'b00111110101010100111011101001111 ;
        3352:  q   <=  32'b10111101100101100111111010011000 ;
        3353:  q   <=  32'b00111111100001100001110011100101 ;
        3354:  q   <=  32'b01000000000000111100010001101000 ;
        3355:  q   <=  32'b00111100110110101010110000000011 ;
        3356:  q   <=  32'b10111110011101100100101111111111 ;
        3357:  q   <=  32'b00111111100001001110110011000001 ;
        3358:  q   <=  32'b10111111000000011101100110000100 ;
        3359:  q   <=  32'b10111111101111011101010110001110 ;
        3360:  q   <=  32'b10111101110110100001011001010101 ;
        3361:  q   <=  32'b00111110011110110010011001111000 ;
        3362:  q   <=  32'b00111110000101010100101011000100 ;
        3363:  q   <=  32'b10111111100011110001110101101100 ;
        3364:  q   <=  32'b10111111000110001101000100100010 ;
        3365:  q   <=  32'b10111111001011011111001011101111 ;
        3366:  q   <=  32'b00111111011101000111111001110010 ;
        3367:  q   <=  32'b10111110000001011111000010010011 ;
        3368:  q   <=  32'b00111111001001100011111101011010 ;
        3369:  q   <=  32'b00111111000110010011100001001000 ;
        3370:  q   <=  32'b10111110010001010001111011011101 ;
        3371:  q   <=  32'b10111111111111011000101011010001 ;
        3372:  q   <=  32'b00111110101110011101001100001011 ;
        3373:  q   <=  32'b00111111001101000011011000001010 ;
        3374:  q   <=  32'b10111111010000001010101000110001 ;
        3375:  q   <=  32'b10111100100010101001011010000001 ;
        3376:  q   <=  32'b10111110111000100010000111001110 ;
        3377:  q   <=  32'b00111111110110011100010101010110 ;
        3378:  q   <=  32'b10111100111110100110110001001101 ;
        3379:  q   <=  32'b00111110010100001100111111010000 ;
        3380:  q   <=  32'b10111111100001100001111010100101 ;
        3381:  q   <=  32'b10111111001111000100000100111011 ;
        3382:  q   <=  32'b10111111101011011010001111010111 ;
        3383:  q   <=  32'b00111111001110101000010010010101 ;
        3384:  q   <=  32'b00111111000110110111000010011001 ;
        3385:  q   <=  32'b10111111010101000000101010000010 ;
        3386:  q   <=  32'b01000000001110001100111100101001 ;
        3387:  q   <=  32'b00111111011010110100110001110101 ;
        3388:  q   <=  32'b00111110110011111100001110010100 ;
        3389:  q   <=  32'b00111111111101010100010110000011 ;
        3390:  q   <=  32'b11000000000111010010100111111100 ;
        3391:  q   <=  32'b10111101101110100111111101110100 ;
        3392:  q   <=  32'b10111100110010100010110111001110 ;
        3393:  q   <=  32'b00111110010011001011110000001000 ;
        3394:  q   <=  32'b10111111100001001110011101111110 ;
        3395:  q   <=  32'b00111111000001111000010010010101 ;
        3396:  q   <=  32'b11000000000011011110010101000110 ;
        3397:  q   <=  32'b00111101110110111111110100011111 ;
        3398:  q   <=  32'b00111110111000001011100010111100 ;
        3399:  q   <=  32'b10111101001001111110100010110100 ;
        3400:  q   <=  32'b00111110101110101000011010111011 ;
        3401:  q   <=  32'b10111111010000111000000110101111 ;
        3402:  q   <=  32'b00111111000011001010110110011011 ;
        3403:  q   <=  32'b10111110101111111101000010000000 ;
        3404:  q   <=  32'b10111111110101000101111101010001 ;
        3405:  q   <=  32'b10111110100111101101011001001000 ;
        3406:  q   <=  32'b10111111000111101011010010010110 ;
        3407:  q   <=  32'b10111111100000110010010111001101 ;
        3408:  q   <=  32'b00111111000000010100011110010101 ;
        3409:  q   <=  32'b00111101001001011100011100100010 ;
        3410:  q   <=  32'b10111110100000100110110000000000 ;
        3411:  q   <=  32'b10111111000011000011100001101011 ;
        3412:  q   <=  32'b00111111110101101001101010100001 ;
        3413:  q   <=  32'b00111111100101100010010011110101 ;
        3414:  q   <=  32'b10111110010000011001100101001010 ;
        3415:  q   <=  32'b00111101101100010100110011111111 ;
        3416:  q   <=  32'b00111111110000011001101110010001 ;
        3417:  q   <=  32'b00111111111001011000100111100101 ;
        3418:  q   <=  32'b00111111100011010010001010101011 ;
        3419:  q   <=  32'b10111110101001101101010101111010 ;
        3420:  q   <=  32'b10111111000101010011001101011011 ;
        3421:  q   <=  32'b00111111010000000110100000000101 ;
        3422:  q   <=  32'b10111111010111010001110110110001 ;
        3423:  q   <=  32'b10111111100010010001001001110011 ;
        3424:  q   <=  32'b10111110101101011110000110011001 ;
        3425:  q   <=  32'b00111111011101001011010010000110 ;
        3426:  q   <=  32'b00111110001000110001101010111010 ;
        3427:  q   <=  32'b00111110011110101101001000000110 ;
        3428:  q   <=  32'b00111111100011111111011111001100 ;
        3429:  q   <=  32'b00111110011100000100001001001101 ;
        3430:  q   <=  32'b10111111100100011011110001101010 ;
        3431:  q   <=  32'b00111111010101111001001101110010 ;
        3432:  q   <=  32'b00111110111100111110001100010011 ;
        3433:  q   <=  32'b10111101101101010000010110100111 ;
        3434:  q   <=  32'b10111110110100110111100101100111 ;
        3435:  q   <=  32'b10111111000010110110100111001111 ;
        3436:  q   <=  32'b10111100110001001010100110101011 ;
        3437:  q   <=  32'b10111111010011001110111001110110 ;
        3438:  q   <=  32'b10111111000000110001111011101000 ;
        3439:  q   <=  32'b10111111101111100100101101100000 ;
        3440:  q   <=  32'b10111111000001001100010110110111 ;
        3441:  q   <=  32'b10111111001100010111011101110101 ;
        3442:  q   <=  32'b00111111000100111110000011111100 ;
        3443:  q   <=  32'b00111111101110100011110001011011 ;
        3444:  q   <=  32'b00111111100001001000101011000100 ;
        3445:  q   <=  32'b00111111100001011111111001001111 ;
        3446:  q   <=  32'b00111111001011010001110000100010 ;
        3447:  q   <=  32'b00111111000010111110110110011111 ;
        3448:  q   <=  32'b00111111001111111111111101000001 ;
        3449:  q   <=  32'b10111111001110101101011010111010 ;
        3450:  q   <=  32'b00111111010101010100110011000001 ;
        3451:  q   <=  32'b10111111100110010110101000011001 ;
        3452:  q   <=  32'b00111111000111100110011111110000 ;
        3453:  q   <=  32'b10111111010101010001100011111110 ;
        3454:  q   <=  32'b10111111011110000111001001011001 ;
        3455:  q   <=  32'b10111110111010000011001010010001 ;
        3456:  q   <=  32'b10111111101001101011111100011110 ;
        3457:  q   <=  32'b00111100100000101101110110010100 ;
        3458:  q   <=  32'b00111111100011100010101000010100 ;
        3459:  q   <=  32'b10111110011111110101101111011110 ;
        3460:  q   <=  32'b00111110111111011100110010011010 ;
        3461:  q   <=  32'b00111110001001011110110100101000 ;
        3462:  q   <=  32'b00111111100110110001110011110011 ;
        3463:  q   <=  32'b10111110001000100001110101111010 ;
        3464:  q   <=  32'b00111110100101100000000001001100 ;
        3465:  q   <=  32'b01000000000111011110111100001000 ;
        3466:  q   <=  32'b00111111100100101011011111001001 ;
        3467:  q   <=  32'b10111111011011110001000001010111 ;
        3468:  q   <=  32'b00111111100011110101010101011000 ;
        3469:  q   <=  32'b10111111011011001001101000011111 ;
        3470:  q   <=  32'b00111100001000100101000011001101 ;
        3471:  q   <=  32'b00111110100101000010011111100100 ;
        3472:  q   <=  32'b00111111010111101011100010000101 ;
        3473:  q   <=  32'b10111110110010110110010111100101 ;
        3474:  q   <=  32'b00111111000010011011000100001100 ;
        3475:  q   <=  32'b00111111111000101000011010111011 ;
        3476:  q   <=  32'b10111111111100111110011011101110 ;
        3477:  q   <=  32'b10111111100010011101001011100001 ;
        3478:  q   <=  32'b00111111100110001111001111010010 ;
        3479:  q   <=  32'b10111110100101101000000001101001 ;
        3480:  q   <=  32'b10111101000111000110000001010101 ;
        3481:  q   <=  32'b00111111011011001000011011111001 ;
        3482:  q   <=  32'b01000000000011100100011010100010 ;
        3483:  q   <=  32'b10111111101001101010010010000010 ;
        3484:  q   <=  32'b10111111011010001011001110011111 ;
        3485:  q   <=  32'b10111101100111101011100001101000 ;
        3486:  q   <=  32'b00111010000001011100111110001010 ;
        3487:  q   <=  32'b00111101110110101101011100000110 ;
        3488:  q   <=  32'b10111110100111111111101101011001 ;
        3489:  q   <=  32'b00111111100111000001110101100001 ;
        3490:  q   <=  32'b10111111011010001101100100000011 ;
        3491:  q   <=  32'b00111110010100001101111101000000 ;
        3492:  q   <=  32'b00111111011111010110000000010110 ;
        3493:  q   <=  32'b00111110110000000001101000101000 ;
        3494:  q   <=  32'b10111111000111110100001110101001 ;
        3495:  q   <=  32'b00111101111101101110010110001001 ;
        3496:  q   <=  32'b10111110101000101000000110111011 ;
        3497:  q   <=  32'b10111111000110011000010011100001 ;
        3498:  q   <=  32'b00111111101011010011010000100101 ;
        3499:  q   <=  32'b10111110010010100110100101100011 ;
        3500:  q   <=  32'b10111111000100111111011111101111 ;
        3501:  q   <=  32'b10111111010000011000011100110111 ;
        3502:  q   <=  32'b00111101111110000011011100100101 ;
        3503:  q   <=  32'b10111111101111110111011110111010 ;
        3504:  q   <=  32'b10111111110100101011010101010101 ;
        3505:  q   <=  32'b00111110010001011000011011101011 ;
        3506:  q   <=  32'b10111111101001010001011100101011 ;
        3507:  q   <=  32'b10111110110011001011100100000000 ;
        3508:  q   <=  32'b00111111010001101000000011010000 ;
        3509:  q   <=  32'b00111111011011000001001000000101 ;
        3510:  q   <=  32'b00111111110001011011001101011001 ;
        3511:  q   <=  32'b10111111100000010011100101010110 ;
        3512:  q   <=  32'b00111111010110110101000100011011 ;
        3513:  q   <=  32'b00111110101001101000101111110101 ;
        3514:  q   <=  32'b00111111101000000100111111101001 ;
        3515:  q   <=  32'b00111110011000010111000101000000 ;
        3516:  q   <=  32'b00111111010100001011000010111010 ;
        3517:  q   <=  32'b00111111100100011101100010010110 ;
        3518:  q   <=  32'b10111110110100101100101111000111 ;
        3519:  q   <=  32'b10111110111011000001000010111001 ;
        3520:  q   <=  32'b10111111101010100001111001000011 ;
        3521:  q   <=  32'b10111101101100110011001101001011 ;
        3522:  q   <=  32'b00111110101101011111110100000100 ;
        3523:  q   <=  32'b10111111001111100011111001010110 ;
        3524:  q   <=  32'b00111101100100111000010011010010 ;
        3525:  q   <=  32'b10111110101101100111101010000000 ;
        3526:  q   <=  32'b10111110110111010000011010110100 ;
        3527:  q   <=  32'b00111111010001111000001000001101 ;
        3528:  q   <=  32'b00111111010100001111101010100101 ;
        3529:  q   <=  32'b00111111100100101111101110100000 ;
        3530:  q   <=  32'b10111111100010101101111111110111 ;
        3531:  q   <=  32'b10111110000010110110001110100011 ;
        3532:  q   <=  32'b00111111001001111011010000010111 ;
        3533:  q   <=  32'b10111111101001011001000000100001 ;
        3534:  q   <=  32'b00111111111101101001111101101010 ;
        3535:  q   <=  32'b00111110011011101101100110001011 ;
        3536:  q   <=  32'b10111111000010111000011010010101 ;
        3537:  q   <=  32'b00111111100001000011001100110011 ;
        3538:  q   <=  32'b00111110110000010001100000001010 ;
        3539:  q   <=  32'b00111101110111111100000101000010 ;
        3540:  q   <=  32'b10111111001011100010000011010001 ;
        3541:  q   <=  32'b10111111111000011111100001100000 ;
        3542:  q   <=  32'b10111111011101101010110001011111 ;
        3543:  q   <=  32'b10111111001001010100100000101110 ;
        3544:  q   <=  32'b00111110111001111011000110111000 ;
        3545:  q   <=  32'b00111111000111010100111111000001 ;
        3546:  q   <=  32'b10111111010010010000100101110110 ;
        3547:  q   <=  32'b00111111010101000000001101011010 ;
        3548:  q   <=  32'b00111111001010101101101111010111 ;
        3549:  q   <=  32'b10111110000000001000001101001101 ;
        3550:  q   <=  32'b10111111011100111000001110111100 ;
        3551:  q   <=  32'b00111111011001000101110010111011 ;
        3552:  q   <=  32'b10111110000001001101010110111011 ;
        3553:  q   <=  32'b10111111100000011011100111100001 ;
        3554:  q   <=  32'b00111110100000010010101111000011 ;
        3555:  q   <=  32'b00111111000001100000100110110000 ;
        3556:  q   <=  32'b10111111101110110001011010101110 ;
        3557:  q   <=  32'b00111111111011101110011001100000 ;
        3558:  q   <=  32'b11000000000010011000101000010001 ;
        3559:  q   <=  32'b10111111110100010100111101101111 ;
        3560:  q   <=  32'b00111111100111001010110010101000 ;
        3561:  q   <=  32'b00111110101001100111110100110101 ;
        3562:  q   <=  32'b10111110110110111001101001111101 ;
        3563:  q   <=  32'b00111100001111011111110110000101 ;
        3564:  q   <=  32'b00111111001110110011011110101111 ;
        3565:  q   <=  32'b10111111010111100011011010111101 ;
        3566:  q   <=  32'b00111111011011011001101111011101 ;
        3567:  q   <=  32'b00111111001100101000001101011001 ;
        3568:  q   <=  32'b10111101001110001110111110010001 ;
        3569:  q   <=  32'b00111110010000111100110011011010 ;
        3570:  q   <=  32'b10111111001000001111011010011011 ;
        3571:  q   <=  32'b10111111010110110100101100000000 ;
        3572:  q   <=  32'b10111110110001110000010101011011 ;
        3573:  q   <=  32'b00111111100000111010011000101010 ;
        3574:  q   <=  32'b10111110011101010111100100111110 ;
        3575:  q   <=  32'b10111110111001110011101100011001 ;
        3576:  q   <=  32'b10111111011110101011000101000001 ;
        3577:  q   <=  32'b10111111100100010001010011001100 ;
        3578:  q   <=  32'b00111100101101010011011011011111 ;
        3579:  q   <=  32'b00111111100001010010011010010001 ;
        3580:  q   <=  32'b00111111100111011010000101000101 ;
        3581:  q   <=  32'b00111111000011110110011111101011 ;
        3582:  q   <=  32'b10111110100111100011101001010001 ;
        3583:  q   <=  32'b10111110101111000011011010011010 ;
        3584:  q   <=  32'b00111110101110110011010001001011 ;
        3585:  q   <=  32'b00111111011011111111101111111011 ;
        3586:  q   <=  32'b00111111011110010110100000001001 ;
        3587:  q   <=  32'b11000000000001111001110001110011 ;
        3588:  q   <=  32'b10111101001111100101000111010000 ;
        3589:  q   <=  32'b10111111011101110111111011110100 ;
        3590:  q   <=  32'b10111110111100010100011110001101 ;
        3591:  q   <=  32'b00111111110111100001101111101110 ;
        3592:  q   <=  32'b10111111010001110000110000110110 ;
        3593:  q   <=  32'b10111111110101111000011010101100 ;
        3594:  q   <=  32'b00111110001101010100011010010111 ;
        3595:  q   <=  32'b10111101111111101110111000010100 ;
        3596:  q   <=  32'b10111110110101001100001110011011 ;
        3597:  q   <=  32'b00111111011000010010010000101101 ;
        3598:  q   <=  32'b00111111000100001110110111000101 ;
        3599:  q   <=  32'b00111110110000000111100000110001 ;
        3600:  q   <=  32'b10111110100011011100110011100100 ;
        3601:  q   <=  32'b00111110101100110100000000011101 ;
        3602:  q   <=  32'b10111110100101010010011000110110 ;
        3603:  q   <=  32'b00111110001111101000101100111111 ;
        3604:  q   <=  32'b00111111000100111001110000000101 ;
        3605:  q   <=  32'b00111110101011011110011110001110 ;
        3606:  q   <=  32'b10111111001011000011111001100101 ;
        3607:  q   <=  32'b10111111000010010111100110111010 ;
        3608:  q   <=  32'b10111111100001010010001111100011 ;
        3609:  q   <=  32'b00111111011111110100111000000110 ;
        3610:  q   <=  32'b10111100110101010110111100010111 ;
        3611:  q   <=  32'b10111111001010000011000100011001 ;
        3612:  q   <=  32'b00111111001011011000000010111100 ;
        3613:  q   <=  32'b10111111000000101100011000000110 ;
        3614:  q   <=  32'b00111110111001000101101010110111 ;
        3615:  q   <=  32'b00111111110000100010000100010101 ;
        3616:  q   <=  32'b00111111011100000001000011001011 ;
        3617:  q   <=  32'b10111110001001000000000110101111 ;
        3618:  q   <=  32'b10111101111010010010001111110101 ;
        3619:  q   <=  32'b00111111111101111111001111000000 ;
        3620:  q   <=  32'b10111110001011101110010111100001 ;
        3621:  q   <=  32'b00111110100110100011001011000011 ;
        3622:  q   <=  32'b00111110101001101110011111111101 ;
        3623:  q   <=  32'b00111111011011001100001000011000 ;
        3624:  q   <=  32'b00111110010111000111010101001101 ;
        3625:  q   <=  32'b00111110101110111000010100000111 ;
        3626:  q   <=  32'b00111110101001001111000011110110 ;
        3627:  q   <=  32'b01000000001011000001100010100010 ;
        3628:  q   <=  32'b00111111011000000100011000001100 ;
        3629:  q   <=  32'b10111111011000000110000110100110 ;
        3630:  q   <=  32'b10111111100110111101010101001101 ;
        3631:  q   <=  32'b10111111110011101011001100010001 ;
        3632:  q   <=  32'b00111111111010111000011111000001 ;
        3633:  q   <=  32'b10111111010100011010010100011110 ;
        3634:  q   <=  32'b00111111011111011111110010011000 ;
        3635:  q   <=  32'b00111111000010001010100001001000 ;
        3636:  q   <=  32'b10111111110000110110101111001011 ;
        3637:  q   <=  32'b01000000000000010111011010000110 ;
        3638:  q   <=  32'b00111111000011010110001101000100 ;
        3639:  q   <=  32'b00111111111010001111101001101101 ;
        3640:  q   <=  32'b00111110101011110110111100011001 ;
        3641:  q   <=  32'b00111110001101111101111011110111 ;
        3642:  q   <=  32'b10111111100000100111100100000101 ;
        3643:  q   <=  32'b00111101000110100000000111100101 ;
        3644:  q   <=  32'b00111110000011000110101000001101 ;
        3645:  q   <=  32'b10111111110000101011000111010111 ;
        3646:  q   <=  32'b10111100100110101111101011011111 ;
        3647:  q   <=  32'b00111110001001110010101000100011 ;
        3648:  q   <=  32'b10111111001110001001110101010100 ;
        3649:  q   <=  32'b00111110110100100011101010011010 ;
        3650:  q   <=  32'b10111111100110110011011101111110 ;
        3651:  q   <=  32'b10111111000100101110000011101110 ;
        3652:  q   <=  32'b00111101110101111101011111011100 ;
        3653:  q   <=  32'b10111111000110101110011110010011 ;
        3654:  q   <=  32'b00111110110101111111010101110110 ;
        3655:  q   <=  32'b10111110101110011100001000011000 ;
        3656:  q   <=  32'b10111111010111111100011000000011 ;
        3657:  q   <=  32'b00111111011011100111110011101111 ;
        3658:  q   <=  32'b00111111000110011001110001011011 ;
        3659:  q   <=  32'b00111111000100100100010010110001 ;
        3660:  q   <=  32'b00111111001011110110001101100001 ;
        3661:  q   <=  32'b00111111100000010011010010110001 ;
        3662:  q   <=  32'b00111111011111011010100110110100 ;
        3663:  q   <=  32'b00111101000010011111111100010101 ;
        3664:  q   <=  32'b10111110111001101000100111001011 ;
        3665:  q   <=  32'b10111101111000101001111111000010 ;
        3666:  q   <=  32'b00111111100111100111001000100111 ;
        3667:  q   <=  32'b10111111100110010101001101111010 ;
        3668:  q   <=  32'b10111111000100000111110000011110 ;
        3669:  q   <=  32'b00111111100001011000101100100010 ;
        3670:  q   <=  32'b00111111010110001001001110010001 ;
        3671:  q   <=  32'b10111110111111011011011011101011 ;
        3672:  q   <=  32'b10111110010100111100100000000101 ;
        3673:  q   <=  32'b10111110000111111000100100000111 ;
        3674:  q   <=  32'b10111110100011010000000011111001 ;
        3675:  q   <=  32'b11000000000111000101111000110001 ;
        3676:  q   <=  32'b10111110110110101100101000001111 ;
        3677:  q   <=  32'b00111110100111100011110100101001 ;
        3678:  q   <=  32'b01000000000111001110011010011011 ;
        3679:  q   <=  32'b10111111101110110011011101100100 ;
        3680:  q   <=  32'b10111111001000101011001011011001 ;
        3681:  q   <=  32'b10111110110001010101110010110010 ;
        3682:  q   <=  32'b10111111011100010011100100011001 ;
        3683:  q   <=  32'b10111111001011000111110001100100 ;
        3684:  q   <=  32'b10111111111101100100110110011111 ;
        3685:  q   <=  32'b10111101111001100011101100110111 ;
        3686:  q   <=  32'b10111111000001001011110100001001 ;
        3687:  q   <=  32'b00111111000010001111010010011101 ;
        3688:  q   <=  32'b00111101011010110010010010001001 ;
        3689:  q   <=  32'b00111111100010000110110010110010 ;
        3690:  q   <=  32'b00111111110011110111010001001100 ;
        3691:  q   <=  32'b00111101111110011000111001101110 ;
        3692:  q   <=  32'b10111111100111100111100000011111 ;
        3693:  q   <=  32'b00111110011110011111110000001110 ;
        3694:  q   <=  32'b00111111101100101111101000100000 ;
        3695:  q   <=  32'b10111101110000111000011110000101 ;
        3696:  q   <=  32'b00111110110001100111011001111101 ;
        3697:  q   <=  32'b10111111011101110110000001100100 ;
        3698:  q   <=  32'b00111111110000010010110100000100 ;
        3699:  q   <=  32'b00111110110011101100001011100111 ;
        3700:  q   <=  32'b10111110110110000010001011100110 ;
        3701:  q   <=  32'b10111111110101100100011001101100 ;
        3702:  q   <=  32'b10111111001100000000100010000111 ;
        3703:  q   <=  32'b10111111100000110111101011001111 ;
        3704:  q   <=  32'b10111110111111000011000001111111 ;
        3705:  q   <=  32'b00111110101100011001000011011100 ;
        3706:  q   <=  32'b00111111010101000101000001110001 ;
        3707:  q   <=  32'b00111110000111110101111000100100 ;
        3708:  q   <=  32'b00111101101010110111001000101100 ;
        3709:  q   <=  32'b00111110101111111100110111000101 ;
        3710:  q   <=  32'b01000000001010011100111000010000 ;
        3711:  q   <=  32'b00111110101010100101100101111100 ;
        3712:  q   <=  32'b00111110000100000010011000111010 ;
        3713:  q   <=  32'b00111111110010011111011001111111 ;
        3714:  q   <=  32'b00111101101101110110010011001110 ;
        3715:  q   <=  32'b10111111001011000100100010101001 ;
        3716:  q   <=  32'b00111111011011101001000010010001 ;
        3717:  q   <=  32'b10111110101101110011110101101000 ;
        3718:  q   <=  32'b00111110010011101111001110111100 ;
        3719:  q   <=  32'b00111111011000000101000111110001 ;
        3720:  q   <=  32'b00111111010011101101010110110011 ;
        3721:  q   <=  32'b10111111110011010011101000001011 ;
        3722:  q   <=  32'b11000000000101110010101111011011 ;
        3723:  q   <=  32'b10111111001100111010001010011110 ;
        3724:  q   <=  32'b00111111110100110111000110010001 ;
        3725:  q   <=  32'b00111110011100001011011011101111 ;
        3726:  q   <=  32'b10111110000110110110010100010100 ;
        3727:  q   <=  32'b10111110000111111010000101000011 ;
        3728:  q   <=  32'b00111111100001001110001010010100 ;
        3729:  q   <=  32'b00111110101010010011010100101011 ;
        3730:  q   <=  32'b00111110111100111001110011101101 ;
        3731:  q   <=  32'b11000000000001011100101011001000 ;
        3732:  q   <=  32'b10111110001100100011011000101110 ;
        3733:  q   <=  32'b00111100100111010011000010000100 ;
        3734:  q   <=  32'b10111111010111000010101011000000 ;
        3735:  q   <=  32'b10111100101111000000000001111000 ;
        3736:  q   <=  32'b10111111000110100011000101110110 ;
        3737:  q   <=  32'b00111111010111101011000111100010 ;
        3738:  q   <=  32'b10111111000100100010000011000011 ;
        3739:  q   <=  32'b00111111101001101111111110111100 ;
        3740:  q   <=  32'b10111101001011101010101110110110 ;
        3741:  q   <=  32'b00111111011001010100000110000001 ;
        3742:  q   <=  32'b01000000000100100011101100010100 ;
        3743:  q   <=  32'b00111101100010001101110011001011 ;
        3744:  q   <=  32'b00111111101111110100111010110100 ;
        3745:  q   <=  32'b10111111100010010100011010000010 ;
        3746:  q   <=  32'b00111111111010010110001101011011 ;
        3747:  q   <=  32'b10111111100110101010110111001110 ;
        3748:  q   <=  32'b10111101100001011110110000000111 ;
        3749:  q   <=  32'b10111110101001110101011100010111 ;
        3750:  q   <=  32'b10111111100100110001011101011110 ;
        3751:  q   <=  32'b10111111101001110110110111101001 ;
        3752:  q   <=  32'b00111111001001010111100101011010 ;
        3753:  q   <=  32'b10111111101100011101000101101011 ;
        3754:  q   <=  32'b10111111101010111001101101111100 ;
        3755:  q   <=  32'b00111111100100000111111011100000 ;
        3756:  q   <=  32'b00111010110111100101000010101001 ;
        3757:  q   <=  32'b00111110110000100110010111101101 ;
        3758:  q   <=  32'b10111111011001101011110110101011 ;
        3759:  q   <=  32'b10111110010010011000010001110100 ;
        3760:  q   <=  32'b00111110100111010010011101101111 ;
        3761:  q   <=  32'b00111110001010110111100111000011 ;
        3762:  q   <=  32'b00111111111001001101111111000100 ;
        3763:  q   <=  32'b10111111000111111100001111011110 ;
        3764:  q   <=  32'b10111110000110011000111101011010 ;
        3765:  q   <=  32'b00111111010101010000110000001011 ;
        3766:  q   <=  32'b00111111011100101011011000011001 ;
        3767:  q   <=  32'b10111111111111001010001101101110 ;
        3768:  q   <=  32'b10111110110010001010010001010001 ;
        3769:  q   <=  32'b10111111001011010011110011110010 ;
        3770:  q   <=  32'b10111100100000110011111001110010 ;
        3771:  q   <=  32'b00111111000000111110001001111110 ;
        3772:  q   <=  32'b00111110111000111100000010110110 ;
        3773:  q   <=  32'b00111111100100100000100011110100 ;
        3774:  q   <=  32'b00111110111001010011011001110010 ;
        3775:  q   <=  32'b00111110101000011000000101100010 ;
        3776:  q   <=  32'b00111111011100100001001001001001 ;
        3777:  q   <=  32'b00111110110110110111100110111011 ;
        3778:  q   <=  32'b10111111101010011000110010111000 ;
        3779:  q   <=  32'b00111101111000001110101000011010 ;
        3780:  q   <=  32'b10111111110100111100110111101101 ;
        3781:  q   <=  32'b00111111100011100010101010000001 ;
        3782:  q   <=  32'b11000000000001101110011100110100 ;
        3783:  q   <=  32'b10111111000011001100001000011101 ;
        3784:  q   <=  32'b00111101110000010000101111000110 ;
        3785:  q   <=  32'b10111101000111001000110001011101 ;
        3786:  q   <=  32'b00111111111100010000001111000011 ;
        3787:  q   <=  32'b00111101011000110010101010111110 ;
        3788:  q   <=  32'b10111111000111010010011111100111 ;
        3789:  q   <=  32'b00111111000101100100011010111000 ;
        3790:  q   <=  32'b10111111100110100111010101101111 ;
        3791:  q   <=  32'b00111111000010111001101011001000 ;
        3792:  q   <=  32'b00111110100000000111100111110010 ;
        3793:  q   <=  32'b10111110110010010001011000110010 ;
        3794:  q   <=  32'b10111111000111110011111000100011 ;
        3795:  q   <=  32'b10111111100110000110000110001010 ;
        3796:  q   <=  32'b10111111111100000111000110011000 ;
        3797:  q   <=  32'b10111110110110010001011110100001 ;
        3798:  q   <=  32'b00111111010001101111100101010011 ;
        3799:  q   <=  32'b10111111001101101100001111011010 ;
        3800:  q   <=  32'b00111111110010101101010101111001 ;
        3801:  q   <=  32'b10111111011000110110100001011110 ;
        3802:  q   <=  32'b01000000000010010000001101011001 ;
        3803:  q   <=  32'b10111111001100010011001010010101 ;
        3804:  q   <=  32'b00111101110010110101110001101000 ;
        3805:  q   <=  32'b00111111101101111010110101011111 ;
        3806:  q   <=  32'b00111111100111011110000000010110 ;
        3807:  q   <=  32'b10111111010000011111010011111110 ;
        3808:  q   <=  32'b00111111001111010001001101110101 ;
        3809:  q   <=  32'b10111111100011101010001101100011 ;
        3810:  q   <=  32'b10111111110110100101100111101011 ;
        3811:  q   <=  32'b00111111001010010100000111101111 ;
        3812:  q   <=  32'b10111111110111010110010011101000 ;
        3813:  q   <=  32'b11000000000010001101011000110010 ;
        3814:  q   <=  32'b10111101011101011111010010001010 ;
        3815:  q   <=  32'b00111111101100010101111001010000 ;
        3816:  q   <=  32'b00111111100110111110000101100011 ;
        3817:  q   <=  32'b10111111101111110101110111010011 ;
        3818:  q   <=  32'b00111101000110001011011000101001 ;
        3819:  q   <=  32'b00111111010011011000100011110010 ;
        3820:  q   <=  32'b00111111011110010100111001110111 ;
        3821:  q   <=  32'b00111111110001111100011000100000 ;
        3822:  q   <=  32'b00111111110010110000101000111001 ;
        3823:  q   <=  32'b00111111010110110011011001010100 ;
        3824:  q   <=  32'b10111111101101100101010101110101 ;
        3825:  q   <=  32'b00111101001000101001111011101011 ;
        3826:  q   <=  32'b10111111101100001010000011110001 ;
        3827:  q   <=  32'b00111111100111011101010101000100 ;
        3828:  q   <=  32'b00111111110111101111110001011011 ;
        3829:  q   <=  32'b11000000000000000001100001111110 ;
        3830:  q   <=  32'b00111111010101011110001100100001 ;
        3831:  q   <=  32'b10111110101011111000010111100010 ;
        3832:  q   <=  32'b10111110111101001011011101110010 ;
        3833:  q   <=  32'b10111111011000111001110000100110 ;
        3834:  q   <=  32'b00111111101000011011100000001011 ;
        3835:  q   <=  32'b00111110110001000011001011110001 ;
        3836:  q   <=  32'b10111101111100110111000010111010 ;
        3837:  q   <=  32'b00111110110101011010000101101011 ;
        3838:  q   <=  32'b00111111100000011011000101000000 ;
        3839:  q   <=  32'b10111111010111101001100010110010 ;
        3840:  q   <=  32'b10111111010010110111000000101110 ;
        3841:  q   <=  32'b00111111001100000100000110101111 ;
        3842:  q   <=  32'b00111111110010101111011101010100 ;
        3843:  q   <=  32'b00111111101000000000010111011100 ;
        3844:  q   <=  32'b10111101111011001100000110001000 ;
        3845:  q   <=  32'b10111111101010100111011101101110 ;
        3846:  q   <=  32'b11000000000101011111000010000110 ;
        3847:  q   <=  32'b10111111011011010011001101000001 ;
        3848:  q   <=  32'b00111111100100001001010110101011 ;
        3849:  q   <=  32'b10111111000011001001001110011111 ;
        3850:  q   <=  32'b00111110100100010100010101001000 ;
        3851:  q   <=  32'b00111110010110011110001011010010 ;
        3852:  q   <=  32'b11000000000011001111101000010010 ;
        3853:  q   <=  32'b00111111101000000010001100101001 ;
        3854:  q   <=  32'b01000000000000011001010011000100 ;
        3855:  q   <=  32'b10111101000111110101001000101001 ;
        3856:  q   <=  32'b00111111011111111010001100101101 ;
        3857:  q   <=  32'b10111111010000011110000010011110 ;
        3858:  q   <=  32'b00111111000110001001110011110111 ;
        3859:  q   <=  32'b01000000000001111110001011001001 ;
        3860:  q   <=  32'b00111111101001111110011010011101 ;
        3861:  q   <=  32'b10111111001100110010111101011101 ;
        3862:  q   <=  32'b10111111100000101000001010110000 ;
        3863:  q   <=  32'b00111101010110011000111011100100 ;
        3864:  q   <=  32'b10111110011100101011010100100111 ;
        3865:  q   <=  32'b10111101100000000111101110111001 ;
        3866:  q   <=  32'b00111111101000101011001110110011 ;
        3867:  q   <=  32'b00111110011000100111001000011000 ;
        3868:  q   <=  32'b00111111110101001111111010110110 ;
        3869:  q   <=  32'b10111101001011111111011010110001 ;
        3870:  q   <=  32'b10111110000010000110111011011111 ;
        3871:  q   <=  32'b00111111010010110000111100100100 ;
        3872:  q   <=  32'b00111110110110100100000001100101 ;
        3873:  q   <=  32'b10111110010101101111000010000011 ;
        3874:  q   <=  32'b10111111110010110100100011001011 ;
        3875:  q   <=  32'b10111111100011101110010110001111 ;
        3876:  q   <=  32'b00111111000111011110101000110110 ;
        3877:  q   <=  32'b00111111000010110010000001111001 ;
        3878:  q   <=  32'b10111111101110111110010000000011 ;
        3879:  q   <=  32'b00111101111101011001001010000000 ;
        3880:  q   <=  32'b00111111000001111000001111010111 ;
        3881:  q   <=  32'b10111111100101100110111001100111 ;
        3882:  q   <=  32'b10111111011111111000101100001000 ;
        3883:  q   <=  32'b00111111100110001101011001100000 ;
        3884:  q   <=  32'b10111111111000000111100100101000 ;
        3885:  q   <=  32'b00111110111001001001111101111110 ;
        3886:  q   <=  32'b00111111011110100110001000100010 ;
        3887:  q   <=  32'b10111111111001010100011111101011 ;
        3888:  q   <=  32'b10111110000001010101000001000100 ;
        3889:  q   <=  32'b10111111100101100110111000101101 ;
        3890:  q   <=  32'b00111101101110000011111000001010 ;
        3891:  q   <=  32'b10111110110110000010011000100000 ;
        3892:  q   <=  32'b10111111110100110101000111001010 ;
        3893:  q   <=  32'b00111111000111100011001100110001 ;
        3894:  q   <=  32'b00111111000110001001110111110101 ;
        3895:  q   <=  32'b10111111000111100101000111101000 ;
        3896:  q   <=  32'b00111111000001110010001011010111 ;
        3897:  q   <=  32'b10111111101011000001001010011101 ;
        3898:  q   <=  32'b10111111100111100000110011001010 ;
        3899:  q   <=  32'b10111111100100111010001111101011 ;
        3900:  q   <=  32'b10111101110111111110011101100001 ;
        3901:  q   <=  32'b10111111000001100011000110100000 ;
        3902:  q   <=  32'b00111111111101001010010101101101 ;
        3903:  q   <=  32'b10111101100100011010000000001010 ;
        3904:  q   <=  32'b00111111000011111101010001110001 ;
        3905:  q   <=  32'b00111111000100101111011001011101 ;
        3906:  q   <=  32'b00111110101111100101001111011100 ;
        3907:  q   <=  32'b00111110010001000100101101100110 ;
        3908:  q   <=  32'b00111111100111110011111000101110 ;
        3909:  q   <=  32'b10111111100101010000001100110000 ;
        3910:  q   <=  32'b00111111110100010101000010000100 ;
        3911:  q   <=  32'b00111111001011111011001101001101 ;
        3912:  q   <=  32'b10111111100100110010001001100000 ;
        3913:  q   <=  32'b00111111100011100001100110100010 ;
        3914:  q   <=  32'b00111111100101110101111000111111 ;
        3915:  q   <=  32'b00111111110110101000100110111010 ;
        3916:  q   <=  32'b10111110110101110011001110010101 ;
        3917:  q   <=  32'b00111111110100011101011100100001 ;
        3918:  q   <=  32'b00111110100001101110010101011000 ;
        3919:  q   <=  32'b10111111101110110101001101101001 ;
        3920:  q   <=  32'b10111111010001101011001100100100 ;
        3921:  q   <=  32'b00111111011011011111001011101101 ;
        3922:  q   <=  32'b00111111111001010111111110100011 ;
        3923:  q   <=  32'b10111111100101110111000110000100 ;
        3924:  q   <=  32'b10111101111000111011000000101011 ;
        3925:  q   <=  32'b10111111001010000010000111001101 ;
        3926:  q   <=  32'b00111111111100001001101100100000 ;
        3927:  q   <=  32'b10111111011001010110010110001110 ;
        3928:  q   <=  32'b00111111101010100110111011000111 ;
        3929:  q   <=  32'b10111111000111111110010000000110 ;
        3930:  q   <=  32'b00111111010001101101010001101101 ;
        3931:  q   <=  32'b10111111101010011000000100100101 ;
        3932:  q   <=  32'b00111111110000000000100100010000 ;
        3933:  q   <=  32'b11000000000011001111110001011100 ;
        3934:  q   <=  32'b00111110101001010010000010100101 ;
        3935:  q   <=  32'b00111110110101111000110111100101 ;
        3936:  q   <=  32'b10111111010100100001100101111000 ;
        3937:  q   <=  32'b10111111011101110110100111010111 ;
        3938:  q   <=  32'b00111111000110111111111000111110 ;
        3939:  q   <=  32'b10111111100001001010001010010011 ;
        3940:  q   <=  32'b10111100111001110101001001011110 ;
        3941:  q   <=  32'b11000000001101000111011100001111 ;
        3942:  q   <=  32'b11000000000001010010111111101010 ;
        3943:  q   <=  32'b10111101001101110100111100001110 ;
        3944:  q   <=  32'b00111111100011110001100100100110 ;
        3945:  q   <=  32'b10111111110100110010001011101110 ;
        3946:  q   <=  32'b00111111001011011011110100100010 ;
        3947:  q   <=  32'b00111110111111010001011111101111 ;
        3948:  q   <=  32'b10111111000101101010010111100000 ;
        3949:  q   <=  32'b10111100110000111111110110100110 ;
        3950:  q   <=  32'b01000000000011000011111001111000 ;
        3951:  q   <=  32'b10111111101100110100011000111101 ;
        3952:  q   <=  32'b00111110111101011100111110011001 ;
        3953:  q   <=  32'b00111110010101001000100000101010 ;
        3954:  q   <=  32'b00111110101001001110100001001011 ;
        3955:  q   <=  32'b10111011110000001011000100010000 ;
        3956:  q   <=  32'b00111110100100000001001000111010 ;
        3957:  q   <=  32'b10111110100000001010111110001001 ;
        3958:  q   <=  32'b10111111110110001100001101000111 ;
        3959:  q   <=  32'b10111111000101011000001000010101 ;
        3960:  q   <=  32'b00111110011100000001000111000001 ;
        3961:  q   <=  32'b00111110100001000111111110100000 ;
        3962:  q   <=  32'b00111111000110101000100100111010 ;
        3963:  q   <=  32'b01000000000011100010010001001011 ;
        3964:  q   <=  32'b10111111110100111011101010001101 ;
        3965:  q   <=  32'b00111111001011100010111101100001 ;
        3966:  q   <=  32'b00111110000010110001011011010110 ;
        3967:  q   <=  32'b10111101000110111001100010111011 ;
        3968:  q   <=  32'b10111111001100010111000101110001 ;
        3969:  q   <=  32'b10111110000000101001010111101010 ;
        3970:  q   <=  32'b00111111001011100010110000110001 ;
        3971:  q   <=  32'b00111110110110100011100011001100 ;
        3972:  q   <=  32'b10111111110011011000011010010011 ;
        3973:  q   <=  32'b00111111011001111111110101101101 ;
        3974:  q   <=  32'b00111110011111111000000010100010 ;
        3975:  q   <=  32'b00111111111100100111011000010001 ;
        3976:  q   <=  32'b10111111100011100110001001101100 ;
        3977:  q   <=  32'b10111111001110001101011110111010 ;
        3978:  q   <=  32'b10111111111000000100011110101000 ;
        3979:  q   <=  32'b00111011011011001011110010010000 ;
        3980:  q   <=  32'b00111111011111101100000111000110 ;
        3981:  q   <=  32'b10111110111101010011101101111000 ;
        3982:  q   <=  32'b10111111000001001110001111010011 ;
        3983:  q   <=  32'b10111110100101101101110110100100 ;
        3984:  q   <=  32'b10111110001001000110011100110010 ;
        3985:  q   <=  32'b00111111100000110000001010010010 ;
        3986:  q   <=  32'b00111100100000100011010110101101 ;
        3987:  q   <=  32'b10111110111101110001111011010011 ;
        3988:  q   <=  32'b00111111001000100111101000000111 ;
        3989:  q   <=  32'b10111111101011101010010111100111 ;
        3990:  q   <=  32'b00111111000110010011111101111001 ;
        3991:  q   <=  32'b10111110010100110111010000111101 ;
        3992:  q   <=  32'b01000000000010001110101101100000 ;
        3993:  q   <=  32'b10111111001001100001100010101000 ;
        3994:  q   <=  32'b00111110110110001110000100010101 ;
        3995:  q   <=  32'b00111101111100010110001101100011 ;
        3996:  q   <=  32'b10111111100010100101011011110010 ;
        3997:  q   <=  32'b00111111011000000010001010000100 ;
        3998:  q   <=  32'b11000000000011100111101101100110 ;
        3999:  q   <=  32'b10111111111110010001101000101100 ;
        4000:  q   <=  32'b10111111101001111010000011001100;
        default: q <= 0;
    endcase
end
endmodule
