module mem_window_cof (clk, addr, cen, wen, data,q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00111101101000111101011100001010 ;
        2:  q   <=  32'b00111101101001000000010111010001 ;
        3:  q   <=  32'b00111101101001001001001000100100 ;
        4:  q   <=  32'b00111101101001010111101111110011 ;
        5:  q   <=  32'b00111101101001101100001100101001 ;
        6:  q   <=  32'b00111101101010000110011110100011 ;
        7:  q   <=  32'b00111101101010100110100100111000 ;
        8:  q   <=  32'b00111101101011001100011110110111 ;
        9:  q   <=  32'b00111101101011111000001011100001 ;
        10:  q   <=  32'b00111101101100101001101001110010 ;
        11:  q   <=  32'b00111101101101100000111000011011 ;
        12:  q   <=  32'b00111101101110011101110110000100 ;
        13:  q   <=  32'b00111101101111100000100001001101 ;
        14:  q   <=  32'b00111101110000101000111000001100 ;
        15:  q   <=  32'b00111101110001110110111001001101 ;
        16:  q   <=  32'b00111101110011001010100010010100 ;
        17:  q   <=  32'b00111101110100100011110001011110 ;
        18:  q   <=  32'b00111101110110000010100100011011 ;
        19:  q   <=  32'b00111101110111100110111000110101 ;
        20:  q   <=  32'b00111101111001010000101100001110 ;
        21:  q   <=  32'b00111101111010111111111011111100 ;
        22:  q   <=  32'b00111101111100110100100101001111 ;
        23:  q   <=  32'b00111101111110101110100101001110 ;
        24:  q   <=  32'b00111110000000010110111100011011 ;
        25:  q   <=  32'b00111110000001011001001110011111 ;
        26:  q   <=  32'b00111110000010011110000111001001 ;
        27:  q   <=  32'b00111110000011100101100100101100 ;
        28:  q   <=  32'b00111110000100101111100101010111 ;
        29:  q   <=  32'b00111110000101111100000111010100 ;
        30:  q   <=  32'b00111110000111001011001000101000 ;
        31:  q   <=  32'b00111110001000011100100111011000 ;
        32:  q   <=  32'b00111110001001110000100001100000 ;
        33:  q   <=  32'b00111110001011000110110100111100 ;
        34:  q   <=  32'b00111110001100011111011111100011 ;
        35:  q   <=  32'b00111110001101111010011111001000 ;
        36:  q   <=  32'b00111110001111010111110001011010 ;
        37:  q   <=  32'b00111110010000110111010100000101 ;
        38:  q   <=  32'b00111110010010011001000100110001 ;
        39:  q   <=  32'b00111110010011111101000001000011 ;
        40:  q   <=  32'b00111110010101100011000110011100 ;
        41:  q   <=  32'b00111110010111001011010010011010 ;
        42:  q   <=  32'b00111110011000110101100010010111 ;
        43:  q   <=  32'b00111110011010100001110011101011 ;
        44:  q   <=  32'b00111110011100010000000011101000 ;
        45:  q   <=  32'b00111110011110000000001111100001 ;
        46:  q   <=  32'b00111110011111110010010100100011 ;
        47:  q   <=  32'b00111110100000110011000111111100 ;
        48:  q   <=  32'b00111110100001101101111111010101 ;
        49:  q   <=  32'b00111110100010101001101110111101 ;
        50:  q   <=  32'b00111110100011100110010101010111 ;
        51:  q   <=  32'b00111110100100100011110001000010 ;
        52:  q   <=  32'b00111110100101100010000000011100 ;
        53:  q   <=  32'b00111110100110100001000010000011 ;
        54:  q   <=  32'b00111110100111100000110100010010 ;
        55:  q   <=  32'b00111110101000100001010101100100 ;
        56:  q   <=  32'b00111110101001100010100100010010 ;
        57:  q   <=  32'b00111110101010100100011110110101 ;
        58:  q   <=  32'b00111110101011100111000011100101 ;
        59:  q   <=  32'b00111110101100101010010000110110 ;
        60:  q   <=  32'b00111110101101101110000100111111 ;
        61:  q   <=  32'b00111110101110110010011110010011 ;
        62:  q   <=  32'b00111110101111110111011011000111 ;
        63:  q   <=  32'b00111110110000111100111001101100 ;
        64:  q   <=  32'b00111110110010000010111000010100 ;
        65:  q   <=  32'b00111110110011001001010101010000 ;
        66:  q   <=  32'b00111110110100010000001110101111 ;
        67:  q   <=  32'b00111110110101010111100011000011 ;
        68:  q   <=  32'b00111110110110011111010000010111 ;
        69:  q   <=  32'b00111110110111100111010100111100 ;
        70:  q   <=  32'b00111110111000101111101110111111 ;
        71:  q   <=  32'b00111110111001111000011100101100 ;
        72:  q   <=  32'b00111110111011000001011100001111 ;
        73:  q   <=  32'b00111110111100001010101011110110 ;
        74:  q   <=  32'b00111110111101010100001001101011 ;
        75:  q   <=  32'b00111110111110011101110011111010 ;
        76:  q   <=  32'b00111110111111100111101000101101 ;
        77:  q   <=  32'b00111111000000011000110011001000 ;
        78:  q   <=  32'b00111111000000111101110101010110 ;
        79:  q   <=  32'b00111111000001100010111010000111 ;
        80:  q   <=  32'b00111111000010001000000000011110 ;
        81:  q   <=  32'b00111111000010101101000111100010 ;
        82:  q   <=  32'b00111111000011010010001110010111 ;
        83:  q   <=  32'b00111111000011110111010100000011 ;
        84:  q   <=  32'b00111111000100011100010111101001 ;
        85:  q   <=  32'b00111111000101000001011000010001 ;
        86:  q   <=  32'b00111111000101100110010100111110 ;
        87:  q   <=  32'b00111111000110001011001100110101 ;
        88:  q   <=  32'b00111111000110101111111110111110 ;
        89:  q   <=  32'b00111111000111010100101010011100 ;
        90:  q   <=  32'b00111111000111111001001110010110 ;
        91:  q   <=  32'b00111111001000011101101001110001 ;
        92:  q   <=  32'b00111111001001000001111011110100 ;
        93:  q   <=  32'b00111111001001100110000011100101 ;
        94:  q   <=  32'b00111111001010001010000000001011 ;
        95:  q   <=  32'b00111111001010101101110000101100 ;
        96:  q   <=  32'b00111111001011010001010100001111 ;
        97:  q   <=  32'b00111111001011110100101001111101 ;
        98:  q   <=  32'b00111111001100010111110000111101 ;
        99:  q   <=  32'b00111111001100111010101000011000 ;
        100:  q   <=  32'b00111111001101011101001111010101 ;
        101:  q   <=  32'b00111111001101111111100100111101 ;
        102:  q   <=  32'b00111111001110100001101000011011 ;
        103:  q   <=  32'b00111111001111000011011000111001 ;
        104:  q   <=  32'b00111111001111100100110101011111 ;
        105:  q   <=  32'b00111111010000000101111101011011 ;
        106:  q   <=  32'b00111111010000100110101111110101 ;
        107:  q   <=  32'b00111111010001000111001011111100 ;
        108:  q   <=  32'b00111111010001100111010000111011 ;
        109:  q   <=  32'b00111111010010000110111101111110 ;
        110:  q   <=  32'b00111111010010100110010010010101 ;
        111:  q   <=  32'b00111111010011000101001101001100 ;
        112:  q   <=  32'b00111111010011100011101101110011 ;
        113:  q   <=  32'b00111111010100000001110011011010 ;
        114:  q   <=  32'b00111111010100011111011101010000 ;
        115:  q   <=  32'b00111111010100111100101010100111 ;
        116:  q   <=  32'b00111111010101011001011010110000 ;
        117:  q   <=  32'b00111111010101110101101100111101 ;
        118:  q   <=  32'b00111111010110010001100000100001 ;
        119:  q   <=  32'b00111111010110101100110100110000 ;
        120:  q   <=  32'b00111111010111000111101001000000 ;
        121:  q   <=  32'b00111111010111100001111100100100 ;
        122:  q   <=  32'b00111111010111111011101110110100 ;
        123:  q   <=  32'b00111111011000010100111111000111 ;
        124:  q   <=  32'b00111111011000101101101100110011 ;
        125:  q   <=  32'b00111111011001000101110111010011 ;
        126:  q   <=  32'b00111111011001011101011101111111 ;
        127:  q   <=  32'b00111111011001110100100000010011 ;
        128:  q   <=  32'b00111111011010001010111101101001 ;
        129:  q   <=  32'b00111111011010100000110101011110 ;
        130:  q   <=  32'b00111111011010110110000111001110 ;
        131:  q   <=  32'b00111111011011001010110010011001 ;
        132:  q   <=  32'b00111111011011011110110110011110 ;
        133:  q   <=  32'b00111111011011110010010010111100 ;
        134:  q   <=  32'b00111111011100000101000111010101 ;
        135:  q   <=  32'b00111111011100010111010011001010 ;
        136:  q   <=  32'b00111111011100101000110101111111 ;
        137:  q   <=  32'b00111111011100111001101111011000 ;
        138:  q   <=  32'b00111111011101001001111110111011 ;
        139:  q   <=  32'b00111111011101011001100100001100 ;
        140:  q   <=  32'b00111111011101101000011110110100 ;
        141:  q   <=  32'b00111111011101110110101110011011 ;
        142:  q   <=  32'b00111111011110000100010010101010 ;
        143:  q   <=  32'b00111111011110010001001011001100 ;
        144:  q   <=  32'b00111111011110011101010111101100 ;
        145:  q   <=  32'b00111111011110101000110111110111 ;
        146:  q   <=  32'b00111111011110110011101011011010 ;
        147:  q   <=  32'b00111111011110111101110010000100 ;
        148:  q   <=  32'b00111111011111000111001011100110 ;
        149:  q   <=  32'b00111111011111001111110111110000 ;
        150:  q   <=  32'b00111111011111010111110110010101 ;
        151:  q   <=  32'b00111111011111011111000111001000 ;
        152:  q   <=  32'b00111111011111100101101001111101 ;
        153:  q   <=  32'b00111111011111101011011110101001 ;
        154:  q   <=  32'b00111111011111110000100101000101 ;
        155:  q   <=  32'b00111111011111110100111101000111 ;
        156:  q   <=  32'b00111111011111111000100110101001 ;
        157:  q   <=  32'b00111111011111111011100001100100 ;
        158:  q   <=  32'b00111111011111111101101101110101 ;
        159:  q   <=  32'b00111111011111111111001011010111 ;
        160:  q   <=  32'b00111111011111111111111010001001 ;
        161:  q   <=  32'b00111111011111111111111010001001 ;
        162:  q   <=  32'b00111111011111111111001011010111 ;
        163:  q   <=  32'b00111111011111111101101101110101 ;
        164:  q   <=  32'b00111111011111111011100001100100 ;
        165:  q   <=  32'b00111111011111111000100110101001 ;
        166:  q   <=  32'b00111111011111110100111101000111 ;
        167:  q   <=  32'b00111111011111110000100101000101 ;
        168:  q   <=  32'b00111111011111101011011110101001 ;
        169:  q   <=  32'b00111111011111100101101001111101 ;
        170:  q   <=  32'b00111111011111011111000111001000 ;
        171:  q   <=  32'b00111111011111010111110110010101 ;
        172:  q   <=  32'b00111111011111001111110111110000 ;
        173:  q   <=  32'b00111111011111000111001011100110 ;
        174:  q   <=  32'b00111111011110111101110010000100 ;
        175:  q   <=  32'b00111111011110110011101011011010 ;
        176:  q   <=  32'b00111111011110101000110111110111 ;
        177:  q   <=  32'b00111111011110011101010111101100 ;
        178:  q   <=  32'b00111111011110010001001011001100 ;
        179:  q   <=  32'b00111111011110000100010010101010 ;
        180:  q   <=  32'b00111111011101110110101110011011 ;
        181:  q   <=  32'b00111111011101101000011110110100 ;
        182:  q   <=  32'b00111111011101011001100100001100 ;
        183:  q   <=  32'b00111111011101001001111110111011 ;
        184:  q   <=  32'b00111111011100111001101111011000 ;
        185:  q   <=  32'b00111111011100101000110101111111 ;
        186:  q   <=  32'b00111111011100010111010011001010 ;
        187:  q   <=  32'b00111111011100000101000111010101 ;
        188:  q   <=  32'b00111111011011110010010010111100 ;
        189:  q   <=  32'b00111111011011011110110110011110 ;
        190:  q   <=  32'b00111111011011001010110010011001 ;
        191:  q   <=  32'b00111111011010110110000111001110 ;
        192:  q   <=  32'b00111111011010100000110101011110 ;
        193:  q   <=  32'b00111111011010001010111101101001 ;
        194:  q   <=  32'b00111111011001110100100000010011 ;
        195:  q   <=  32'b00111111011001011101011101111111 ;
        196:  q   <=  32'b00111111011001000101110111010011 ;
        197:  q   <=  32'b00111111011000101101101100110011 ;
        198:  q   <=  32'b00111111011000010100111111000111 ;
        199:  q   <=  32'b00111111010111111011101110110100 ;
        200:  q   <=  32'b00111111010111100001111100100100 ;
        201:  q   <=  32'b00111111010111000111101001000000 ;
        202:  q   <=  32'b00111111010110101100110100110000 ;
        203:  q   <=  32'b00111111010110010001100000100001 ;
        204:  q   <=  32'b00111111010101110101101100111101 ;
        205:  q   <=  32'b00111111010101011001011010110000 ;
        206:  q   <=  32'b00111111010100111100101010100111 ;
        207:  q   <=  32'b00111111010100011111011101010000 ;
        208:  q   <=  32'b00111111010100000001110011011010 ;
        209:  q   <=  32'b00111111010011100011101101110011 ;
        210:  q   <=  32'b00111111010011000101001101001100 ;
        211:  q   <=  32'b00111111010010100110010010010101 ;
        212:  q   <=  32'b00111111010010000110111101111110 ;
        213:  q   <=  32'b00111111010001100111010000111011 ;
        214:  q   <=  32'b00111111010001000111001011111100 ;
        215:  q   <=  32'b00111111010000100110101111110101 ;
        216:  q   <=  32'b00111111010000000101111101011011 ;
        217:  q   <=  32'b00111111001111100100110101011111 ;
        218:  q   <=  32'b00111111001111000011011000111001 ;
        219:  q   <=  32'b00111111001110100001101000011011 ;
        220:  q   <=  32'b00111111001101111111100100111101 ;
        221:  q   <=  32'b00111111001101011101001111010101 ;
        222:  q   <=  32'b00111111001100111010101000011000 ;
        223:  q   <=  32'b00111111001100010111110000111101 ;
        224:  q   <=  32'b00111111001011110100101001111101 ;
        225:  q   <=  32'b00111111001011010001010100001111 ;
        226:  q   <=  32'b00111111001010101101110000101100 ;
        227:  q   <=  32'b00111111001010001010000000001011 ;
        228:  q   <=  32'b00111111001001100110000011100101 ;
        229:  q   <=  32'b00111111001001000001111011110100 ;
        230:  q   <=  32'b00111111001000011101101001110001 ;
        231:  q   <=  32'b00111111000111111001001110010110 ;
        232:  q   <=  32'b00111111000111010100101010011100 ;
        233:  q   <=  32'b00111111000110101111111110111110 ;
        234:  q   <=  32'b00111111000110001011001100110101 ;
        235:  q   <=  32'b00111111000101100110010100111110 ;
        236:  q   <=  32'b00111111000101000001011000010001 ;
        237:  q   <=  32'b00111111000100011100010111101001 ;
        238:  q   <=  32'b00111111000011110111010100000011 ;
        239:  q   <=  32'b00111111000011010010001110010111 ;
        240:  q   <=  32'b00111111000010101101000111100010 ;
        241:  q   <=  32'b00111111000010001000000000011110 ;
        242:  q   <=  32'b00111111000001100010111010000111 ;
        243:  q   <=  32'b00111111000000111101110101010110 ;
        244:  q   <=  32'b00111111000000011000110011001000 ;
        245:  q   <=  32'b00111110111111100111101000101101 ;
        246:  q   <=  32'b00111110111110011101110011111010 ;
        247:  q   <=  32'b00111110111101010100001001101011 ;
        248:  q   <=  32'b00111110111100001010101011110110 ;
        249:  q   <=  32'b00111110111011000001011100001111 ;
        250:  q   <=  32'b00111110111001111000011100101100 ;
        251:  q   <=  32'b00111110111000101111101110111111 ;
        252:  q   <=  32'b00111110110111100111010100111100 ;
        253:  q   <=  32'b00111110110110011111010000010111 ;
        254:  q   <=  32'b00111110110101010111100011000011 ;
        255:  q   <=  32'b00111110110100010000001110101111 ;
        256:  q   <=  32'b00111110110011001001010101010000 ;
        257:  q   <=  32'b00111110110010000010111000010100 ;
        258:  q   <=  32'b00111110110000111100111001101100 ;
        259:  q   <=  32'b00111110101111110111011011000111 ;
        260:  q   <=  32'b00111110101110110010011110010011 ;
        261:  q   <=  32'b00111110101101101110000100111111 ;
        262:  q   <=  32'b00111110101100101010010000110110 ;
        263:  q   <=  32'b00111110101011100111000011100101 ;
        264:  q   <=  32'b00111110101010100100011110110101 ;
        265:  q   <=  32'b00111110101001100010100100010010 ;
        266:  q   <=  32'b00111110101000100001010101100100 ;
        267:  q   <=  32'b00111110100111100000110100010010 ;
        268:  q   <=  32'b00111110100110100001000010000011 ;
        269:  q   <=  32'b00111110100101100010000000011100 ;
        270:  q   <=  32'b00111110100100100011110001000010 ;
        271:  q   <=  32'b00111110100011100110010101010111 ;
        272:  q   <=  32'b00111110100010101001101110111101 ;
        273:  q   <=  32'b00111110100001101101111111010101 ;
        274:  q   <=  32'b00111110100000110011000111111100 ;
        275:  q   <=  32'b00111110011111110010010100100011 ;
        276:  q   <=  32'b00111110011110000000001111100001 ;
        277:  q   <=  32'b00111110011100010000000011101000 ;
        278:  q   <=  32'b00111110011010100001110011101011 ;
        279:  q   <=  32'b00111110011000110101100010010111 ;
        280:  q   <=  32'b00111110010111001011010010011010 ;
        281:  q   <=  32'b00111110010101100011000110011100 ;
        282:  q   <=  32'b00111110010011111101000001000011 ;
        283:  q   <=  32'b00111110010010011001000100110001 ;
        284:  q   <=  32'b00111110010000110111010100000101 ;
        285:  q   <=  32'b00111110001111010111110001011010 ;
        286:  q   <=  32'b00111110001101111010011111001000 ;
        287:  q   <=  32'b00111110001100011111011111100011 ;
        288:  q   <=  32'b00111110001011000110110100111100 ;
        289:  q   <=  32'b00111110001001110000100001100000 ;
        290:  q   <=  32'b00111110001000011100100111011000 ;
        291:  q   <=  32'b00111110000111001011001000101000 ;
        292:  q   <=  32'b00111110000101111100000111010100 ;
        293:  q   <=  32'b00111110000100101111100101010111 ;
        294:  q   <=  32'b00111110000011100101100100101100 ;
        295:  q   <=  32'b00111110000010011110000111001001 ;
        296:  q   <=  32'b00111110000001011001001110011111 ;
        297:  q   <=  32'b00111110000000010110111100011011 ;
        298:  q   <=  32'b00111101111110101110100101001110 ;
        299:  q   <=  32'b00111101111100110100100101001111 ;
        300:  q   <=  32'b00111101111010111111111011111100 ;
        301:  q   <=  32'b00111101111001010000101100001110 ;
        302:  q   <=  32'b00111101110111100110111000110101 ;
        303:  q   <=  32'b00111101110110000010100100011011 ;
        304:  q   <=  32'b00111101110100100011110001011110 ;
        305:  q   <=  32'b00111101110011001010100010010100 ;
        306:  q   <=  32'b00111101110001110110111001001101 ;
        307:  q   <=  32'b00111101110000101000111000001100 ;
        308:  q   <=  32'b00111101101111100000100001001101 ;
        309:  q   <=  32'b00111101101110011101110110000100 ;
        310:  q   <=  32'b00111101101101100000111000011011 ;
        311:  q   <=  32'b00111101101100101001101001110010 ;
        312:  q   <=  32'b00111101101011111000001011100001 ;
        313:  q   <=  32'b00111101101011001100011110110111 ;
        314:  q   <=  32'b00111101101010100110100100111000 ;
        315:  q   <=  32'b00111101101010000110011110100011 ;
        316:  q   <=  32'b00111101101001101100001100101001 ;
        317:  q   <=  32'b00111101101001010111101111110011 ;
        318:  q   <=  32'b00111101101001001001001000100100 ;
        319:  q   <=  32'b00111101101001000000010111010001 ;
        320:  q   <=  32'b00111101101000111101011100001010;
        default: q <= 0;
    endcase
end
endmodule
