module mem_mel_cof_3 (clk, addr, cen, wen, data, q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;// Note
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        0:  q   <=  32'b00000000000000000000000000000000 ;
        1:  q   <=  32'b00000000000000000000000000000000 ;
        2:  q   <=  32'b00000000000000000000000000000000 ;
        3:  q   <=  32'b00000000000000000000000000000000 ;
        4:  q   <=  32'b00000000000000000000000000000000 ;
        5:  q   <=  32'b00000000000000000000000000000000 ;
        6:  q   <=  32'b00000000000000000000000000000000 ;
        7:  q   <=  32'b00000000000000000000000000000000 ;
        8:  q   <=  32'b00000000000000000000000000000000 ;
        9:  q   <=  32'b00000000000000000000000000000000 ;
        10:  q   <=  32'b00000000000000000000000000000000 ;
        11:  q   <=  32'b00000000000000000000000000000000 ;
        12:  q   <=  32'b00000000000000000000000000000000 ;
        13:  q   <=  32'b00000000000000000000000000000000 ;
        14:  q   <=  32'b00000000000000000000000000000000 ;
        15:  q   <=  32'b00000000000000000000000000000000 ;
        16:  q   <=  32'b00000000000000000000000000000000 ;
        17:  q   <=  32'b00000000000000000000000000000000 ;
        18:  q   <=  32'b00000000000000000000000000000000 ;
        19:  q   <=  32'b00000000000000000000000000000000 ;
        20:  q   <=  32'b00000000000000000000000000000000 ;
        21:  q   <=  32'b00000000000000000000000000000000 ;
        22:  q   <=  32'b00000000000000000000000000000000 ;
        23:  q   <=  32'b00000000000000000000000000000000 ;
        24:  q   <=  32'b00000000000000000000000000000000 ;
        25:  q   <=  32'b00000000000000000000000000000000 ;
        26:  q   <=  32'b00000000000000000000000000000000 ;
        27:  q   <=  32'b00000000000000000000000000000000 ;
        28:  q   <=  32'b00000000000000000000000000000000 ;
        29:  q   <=  32'b00000000000000000000000000000000 ;
        30:  q   <=  32'b00000000000000000000000000000000 ;
        31:  q   <=  32'b00000000000000000000000000000000 ;
        32:  q   <=  32'b00000000000000000000000000000000 ;
        33:  q   <=  32'b00000000000000000000000000000000 ;
        34:  q   <=  32'b00000000000000000000000000000000 ;
        35:  q   <=  32'b00000000000000000000000000000000 ;
        36:  q   <=  32'b00000000000000000000000000000000 ;
        37:  q   <=  32'b00000000000000000000000000000000 ;
        38:  q   <=  32'b00000000000000000000000000000000 ;
        39:  q   <=  32'b00000000000000000000000000000000 ;
        40:  q   <=  32'b00000000000000000000000000000000 ;
        41:  q   <=  32'b00000000000000000000000000000000 ;
        42:  q   <=  32'b00000000000000000000000000000000 ;
        43:  q   <=  32'b00000000000000000000000000000000 ;
        44:  q   <=  32'b00000000000000000000000000000000 ;
        45:  q   <=  32'b00000000000000000000000000000000 ;
        46:  q   <=  32'b00000000000000000000000000000000 ;
        47:  q   <=  32'b00000000000000000000000000000000 ;
        48:  q   <=  32'b00000000000000000000000000000000 ;
        49:  q   <=  32'b00000000000000000000000000000000 ;
        50:  q   <=  32'b00000000000000000000000000000000 ;
        51:  q   <=  32'b00000000000000000000000000000000 ;
        52:  q   <=  32'b00000000000000000000000000000000 ;
        53:  q   <=  32'b00000000000000000000000000000000 ;
        54:  q   <=  32'b00000000000000000000000000000000 ;
        55:  q   <=  32'b00000000000000000000000000000000 ;
        56:  q   <=  32'b00000000000000000000000000000000 ;
        57:  q   <=  32'b00000000000000000000000000000000 ;
        58:  q   <=  32'b00000000000000000000000000000000 ;
        59:  q   <=  32'b00000000000000000000000000000000 ;
        60:  q   <=  32'b00000000000000000000000000000000 ;
        61:  q   <=  32'b00000000000000000000000000000000 ;
        62:  q   <=  32'b00000000000000000000000000000000 ;
        63:  q   <=  32'b00000000000000000000000000000000 ;
        64:  q   <=  32'b00000000000000000000000000000000 ;
        65:  q   <=  32'b00000000000000000000000000000000 ;
        66:  q   <=  32'b00000000000000000000000000000000 ;
        67:  q   <=  32'b00000000000000000000000000000000 ;
        68:  q   <=  32'b00000000000000000000000000000000 ;
        69:  q   <=  32'b00000000000000000000000000000000 ;
        70:  q   <=  32'b00000000000000000000000000000000 ;
        71:  q   <=  32'b00000000000000000000000000000000 ;
        72:  q   <=  32'b00000000000000000000000000000000 ;
        73:  q   <=  32'b00000000000000000000000000000000 ;
        74:  q   <=  32'b00000000000000000000000000000000 ;
        75:  q   <=  32'b00000000000000000000000000000000 ;
        76:  q   <=  32'b00000000000000000000000000000000 ;
        77:  q   <=  32'b00000000000000000000000000000000 ;
        78:  q   <=  32'b00000000000000000000000000000000 ;
        79:  q   <=  32'b00000000000000000000000000000000 ;
        80:  q   <=  32'b00000000000000000000000000000000 ;
        81:  q   <=  32'b00000000000000000000000000000000 ;
        82:  q   <=  32'b00000000000000000000000000000000 ;
        83:  q   <=  32'b00000000000000000000000000000000 ;
        84:  q   <=  32'b00000000000000000000000000000000 ;
        85:  q   <=  32'b00000000000000000000000000000000 ;
        86:  q   <=  32'b00000000000000000000000000000000 ;
        87:  q   <=  32'b00000000000000000000000000000000 ;
        88:  q   <=  32'b00000000000000000000000000000000 ;
        89:  q   <=  32'b00000000000000000000000000000000 ;
        90:  q   <=  32'b00000000000000000000000000000000 ;
        91:  q   <=  32'b00000000000000000000000000000000 ;
        92:  q   <=  32'b00000000000000000000000000000000 ;
        93:  q   <=  32'b00000000000000000000000000000000 ;
        94:  q   <=  32'b00000000000000000000000000000000 ;
        95:  q   <=  32'b00000000000000000000000000000000 ;
        96:  q   <=  32'b00000000000000000000000000000000 ;
        97:  q   <=  32'b00000000000000000000000000000000 ;
        98:  q   <=  32'b00000000000000000000000000000000 ;
        99:  q   <=  32'b00000000000000000000000000000000 ;
        100:  q   <=  32'b00000000000000000000000000000000 ;
        101:  q   <=  32'b00000000000000000000000000000000 ;
        102:  q   <=  32'b00000000000000000000000000000000 ;
        103:  q   <=  32'b00000000000000000000000000000000 ;
        104:  q   <=  32'b00000000000000000000000000000000 ;
        105:  q   <=  32'b00000000000000000000000000000000 ;
        106:  q   <=  32'b00000000000000000000000000000000 ;
        107:  q   <=  32'b00000000000000000000000000000000 ;
        108:  q   <=  32'b00000000000000000000000000000000 ;
        109:  q   <=  32'b00000000000000000000000000000000 ;
        110:  q   <=  32'b00000000000000000000000000000000 ;
        111:  q   <=  32'b00000000000000000000000000000000 ;
        112:  q   <=  32'b00000000000000000000000000000000 ;
        113:  q   <=  32'b00000000000000000000000000000000 ;
        114:  q   <=  32'b00000000000000000000000000000000 ;
        115:  q   <=  32'b00000000000000000000000000000000 ;
        116:  q   <=  32'b00000000000000000000000000000000 ;
        117:  q   <=  32'b00000000000000000000000000000000 ;
        118:  q   <=  32'b00000000000000000000000000000000 ;
        119:  q   <=  32'b00000000000000000000000000000000 ;
        120:  q   <=  32'b00000000000000000000000000000000 ;
        121:  q   <=  32'b00000000000000000000000000000000 ;
        122:  q   <=  32'b00000000000000000000000000000000 ;
        123:  q   <=  32'b00000000000000000000000000000000 ;
        124:  q   <=  32'b00000000000000000000000000000000 ;
        125:  q   <=  32'b00000000000000000000000000000000 ;
        126:  q   <=  32'b00000000000000000000000000000000 ;
        127:  q   <=  32'b00000000000000000000000000000000 ;
        128:  q   <=  32'b00000000000000000000000000000000 ;
        129:  q   <=  32'b00000000000000000000000000000000 ;
        130:  q   <=  32'b00111101111111001011000100000100 ;
        131:  q   <=  32'b00111110111111111101011110001011 ;
        132:  q   <=  32'b00111111010111111000000111010011 ;
        133:  q   <=  32'b00111111100111110010110101000001 ;
        134:  q   <=  32'b00111111110011100011110000000011 ;
        135:  q   <=  32'b00111111111111001110111001000001 ;
        136:  q   <=  32'b00111111110101001011101011110011 ;
        137:  q   <=  32'b00111111101001101011111010001111 ;
        138:  q   <=  32'b00111111011100100011011100010101 ;
        139:  q   <=  32'b00111111000101111010000111000101 ;
        140:  q   <=  32'b00111110011101101110110010111101 ;
        141:  q   <=  32'b00000000000000000000000000000000 ;
        142:  q   <=  32'b00000000000000000000000000000000 ;
        143:  q   <=  32'b00000000000000000000000000000000 ;
        144:  q   <=  32'b00000000000000000000000000000000 ;
        145:  q   <=  32'b00000000000000000000000000000000 ;
        146:  q   <=  32'b00000000000000000000000000000000 ;
        147:  q   <=  32'b00000000000000000000000000000000 ;
        148:  q   <=  32'b00000000000000000000000000000000 ;
        149:  q   <=  32'b00000000000000000000000000000000 ;
        150:  q   <=  32'b00000000000000000000000000000000 ;
        151:  q   <=  32'b00000000000000000000000000000000 ;
        152:  q   <=  32'b00000000000000000000000000000000 ;
        153:  q   <=  32'b00000000000000000000000000000000 ;
        154:  q   <=  32'b00000000000000000000000000000000 ;
        155:  q   <=  32'b00000000000000000000000000000000 ;
        156:  q   <=  32'b00000000000000000000000000000000 ;
        157:  q   <=  32'b00000000000000000000000000000000 ;
        158:  q   <=  32'b00000000000000000000000000000000 ;
        159:  q   <=  32'b00000000000000000000000000000000 ;
        160:  q   <=  32'b00000000000000000000000000000000 ;
        161:  q   <=  32'b00000000000000000000000000000000 ;
        162:  q   <=  32'b00000000000000000000000000000000 ;
        163:  q   <=  32'b00000000000000000000000000000000 ;
        164:  q   <=  32'b00000000000000000000000000000000 ;
        165:  q   <=  32'b00000000000000000000000000000000 ;
        166:  q   <=  32'b00000000000000000000000000000000 ;
        167:  q   <=  32'b00000000000000000000000000000000 ;
        168:  q   <=  32'b00000000000000000000000000000000 ;
        169:  q   <=  32'b00000000000000000000000000000000 ;
        170:  q   <=  32'b00000000000000000000000000000000 ;
        171:  q   <=  32'b00000000000000000000000000000000 ;
        172:  q   <=  32'b00000000000000000000000000000000 ;
        173:  q   <=  32'b00000000000000000000000000000000 ;
        174:  q   <=  32'b00000000000000000000000000000000 ;
        175:  q   <=  32'b00000000000000000000000000000000 ;
        176:  q   <=  32'b00000000000000000000000000000000 ;
        177:  q   <=  32'b00000000000000000000000000000000 ;
        178:  q   <=  32'b00000000000000000000000000000000 ;
        179:  q   <=  32'b00000000000000000000000000000000 ;
        180:  q   <=  32'b00000000000000000000000000000000 ;
        181:  q   <=  32'b00000000000000000000000000000000 ;
        182:  q   <=  32'b00000000000000000000000000000000 ;
        183:  q   <=  32'b00000000000000000000000000000000 ;
        184:  q   <=  32'b00000000000000000000000000000000 ;
        185:  q   <=  32'b00000000000000000000000000000000 ;
        186:  q   <=  32'b00000000000000000000000000000000 ;
        187:  q   <=  32'b00000000000000000000000000000000 ;
        188:  q   <=  32'b00000000000000000000000000000000 ;
        189:  q   <=  32'b00000000000000000000000000000000 ;
        190:  q   <=  32'b00000000000000000000000000000000 ;
        191:  q   <=  32'b00000000000000000000000000000000 ;
        192:  q   <=  32'b00000000000000000000000000000000 ;
        193:  q   <=  32'b00000000000000000000000000000000 ;
        194:  q   <=  32'b00000000000000000000000000000000 ;
        195:  q   <=  32'b00000000000000000000000000000000 ;
        196:  q   <=  32'b00000000000000000000000000000000 ;
        197:  q   <=  32'b00000000000000000000000000000000 ;
        198:  q   <=  32'b00000000000000000000000000000000 ;
        199:  q   <=  32'b00000000000000000000000000000000 ;
        200:  q   <=  32'b00000000000000000000000000000000 ;
        201:  q   <=  32'b00000000000000000000000000000000 ;
        202:  q   <=  32'b00000000000000000000000000000000 ;
        203:  q   <=  32'b00000000000000000000000000000000 ;
        204:  q   <=  32'b00000000000000000000000000000000 ;
        205:  q   <=  32'b00000000000000000000000000000000 ;
        206:  q   <=  32'b00000000000000000000000000000000 ;
        207:  q   <=  32'b00000000000000000000000000000000 ;
        208:  q   <=  32'b00000000000000000000000000000000 ;
        209:  q   <=  32'b00000000000000000000000000000000 ;
        210:  q   <=  32'b00000000000000000000000000000000 ;
        211:  q   <=  32'b00000000000000000000000000000000 ;
        212:  q   <=  32'b00000000000000000000000000000000 ;
        213:  q   <=  32'b00000000000000000000000000000000 ;
        214:  q   <=  32'b00000000000000000000000000000000 ;
        215:  q   <=  32'b00000000000000000000000000000000 ;
        216:  q   <=  32'b00000000000000000000000000000000 ;
        217:  q   <=  32'b00000000000000000000000000000000 ;
        218:  q   <=  32'b00000000000000000000000000000000 ;
        219:  q   <=  32'b00000000000000000000000000000000 ;
        220:  q   <=  32'b00000000000000000000000000000000 ;
        221:  q   <=  32'b00000000000000000000000000000000 ;
        222:  q   <=  32'b00000000000000000000000000000000 ;
        223:  q   <=  32'b00000000000000000000000000000000 ;
        224:  q   <=  32'b00000000000000000000000000000000 ;
        225:  q   <=  32'b00000000000000000000000000000000 ;
        226:  q   <=  32'b00000000000000000000000000000000 ;
        227:  q   <=  32'b00000000000000000000000000000000 ;
        228:  q   <=  32'b00000000000000000000000000000000 ;
        229:  q   <=  32'b00000000000000000000000000000000 ;
        230:  q   <=  32'b00000000000000000000000000000000 ;
        231:  q   <=  32'b00000000000000000000000000000000 ;
        232:  q   <=  32'b00000000000000000000000000000000 ;
        233:  q   <=  32'b00000000000000000000000000000000 ;
        234:  q   <=  32'b00000000000000000000000000000000 ;
        235:  q   <=  32'b00000000000000000000000000000000 ;
        236:  q   <=  32'b00000000000000000000000000000000 ;
        237:  q   <=  32'b00000000000000000000000000000000 ;
        238:  q   <=  32'b00000000000000000000000000000000 ;
        239:  q   <=  32'b00000000000000000000000000000000 ;
        240:  q   <=  32'b00000000000000000000000000000000 ;
        241:  q   <=  32'b00000000000000000000000000000000 ;
        242:  q   <=  32'b00000000000000000000000000000000 ;
        243:  q   <=  32'b00000000000000000000000000000000 ;
        244:  q   <=  32'b00000000000000000000000000000000 ;
        245:  q   <=  32'b00000000000000000000000000000000 ;
        246:  q   <=  32'b00000000000000000000000000000000 ;
        247:  q   <=  32'b00000000000000000000000000000000 ;
        248:  q   <=  32'b00000000000000000000000000000000 ;
        249:  q   <=  32'b00000000000000000000000000000000 ;
        250:  q   <=  32'b00000000000000000000000000000000 ;
        251:  q   <=  32'b00000000000000000000000000000000 ;
        252:  q   <=  32'b00000000000000000000000000000000 ;
        253:  q   <=  32'b00000000000000000000000000000000 ;
        254:  q   <=  32'b00000000000000000000000000000000 ;
        255:  q   <=  32'b00000000000000000000000000000000 ;
        256:  q   <=  32'b00000000000000000000000000000000 ;
        257:  q   <=  32'b00000000000000000000000000000000 ;
        258:  q   <=  32'b00000000000000000000000000000000 ;
        259:  q   <=  32'b00000000000000000000000000000000 ;
        260:  q   <=  32'b00000000000000000000000000000000 ;
        261:  q   <=  32'b00000000000000000000000000000000 ;
        262:  q   <=  32'b00000000000000000000000000000000 ;
        263:  q   <=  32'b00000000000000000000000000000000 ;
        264:  q   <=  32'b00000000000000000000000000000000 ;
        265:  q   <=  32'b00000000000000000000000000000000 ;
        266:  q   <=  32'b00000000000000000000000000000000 ;
        267:  q   <=  32'b00000000000000000000000000000000 ;
        268:  q   <=  32'b00000000000000000000000000000000 ;
        269:  q   <=  32'b00000000000000000000000000000000 ;
        270:  q   <=  32'b00000000000000000000000000000000 ;
        271:  q   <=  32'b00000000000000000000000000000000 ;
        272:  q   <=  32'b00000000000000000000000000000000 ;
        273:  q   <=  32'b00000000000000000000000000000000 ;
        274:  q   <=  32'b00000000000000000000000000000000 ;
        275:  q   <=  32'b00000000000000000000000000000000 ;
        276:  q   <=  32'b00000000000000000000000000000000 ;
        277:  q   <=  32'b00000000000000000000000000000000 ;
        278:  q   <=  32'b00000000000000000000000000000000 ;
        279:  q   <=  32'b00000000000000000000000000000000 ;
        280:  q   <=  32'b00000000000000000000000000000000 ;
        281:  q   <=  32'b00000000000000000000000000000000 ;
        282:  q   <=  32'b00000000000000000000000000000000 ;
        283:  q   <=  32'b00000000000000000000000000000000 ;
        284:  q   <=  32'b00000000000000000000000000000000 ;
        285:  q   <=  32'b00000000000000000000000000000000 ;
        286:  q   <=  32'b00000000000000000000000000000000 ;
        287:  q   <=  32'b00000000000000000000000000000000 ;
        288:  q   <=  32'b00000000000000000000000000000000 ;
        289:  q   <=  32'b00000000000000000000000000000000 ;
        290:  q   <=  32'b00000000000000000000000000000000 ;
        291:  q   <=  32'b00000000000000000000000000000000 ;
        292:  q   <=  32'b00000000000000000000000000000000 ;
        293:  q   <=  32'b00000000000000000000000000000000 ;
        294:  q   <=  32'b00000000000000000000000000000000 ;
        295:  q   <=  32'b00000000000000000000000000000000 ;
        296:  q   <=  32'b00000000000000000000000000000000 ;
        297:  q   <=  32'b00000000000000000000000000000000 ;
        298:  q   <=  32'b00000000000000000000000000000000 ;
        299:  q   <=  32'b00000000000000000000000000000000 ;
        300:  q   <=  32'b00000000000000000000000000000000 ;
        301:  q   <=  32'b00000000000000000000000000000000 ;
        302:  q   <=  32'b00000000000000000000000000000000 ;
        303:  q   <=  32'b00000000000000000000000000000000 ;
        304:  q   <=  32'b00000000000000000000000000000000 ;
        305:  q   <=  32'b00000000000000000000000000000000 ;
        306:  q   <=  32'b00000000000000000000000000000000 ;
        307:  q   <=  32'b00000000000000000000000000000000 ;
        308:  q   <=  32'b00000000000000000000000000000000 ;
        309:  q   <=  32'b00000000000000000000000000000000 ;
        310:  q   <=  32'b00000000000000000000000000000000 ;
        311:  q   <=  32'b00000000000000000000000000000000 ;
        312:  q   <=  32'b00000000000000000000000000000000 ;
        313:  q   <=  32'b00000000000000000000000000000000 ;
        314:  q   <=  32'b00000000000000000000000000000000 ;
        315:  q   <=  32'b00000000000000000000000000000000 ;
        316:  q   <=  32'b00000000000000000000000000000000 ;
        317:  q   <=  32'b00000000000000000000000000000000 ;
        318:  q   <=  32'b00000000000000000000000000000000 ;
        319:  q   <=  32'b00000000000000000000000000000000 ;
        320:  q   <=  32'b00000000000000000000000000000000 ;
        321:  q   <=  32'b00000000000000000000000000000000 ;
        322:  q   <=  32'b00000000000000000000000000000000 ;
        323:  q   <=  32'b00000000000000000000000000000000 ;
        324:  q   <=  32'b00000000000000000000000000000000 ;
        325:  q   <=  32'b00000000000000000000000000000000 ;
        326:  q   <=  32'b00000000000000000000000000000000 ;
        327:  q   <=  32'b00000000000000000000000000000000 ;
        328:  q   <=  32'b00000000000000000000000000000000 ;
        329:  q   <=  32'b00000000000000000000000000000000 ;
        330:  q   <=  32'b00000000000000000000000000000000 ;
        331:  q   <=  32'b00000000000000000000000000000000 ;
        332:  q   <=  32'b00000000000000000000000000000000 ;
        333:  q   <=  32'b00000000000000000000000000000000 ;
        334:  q   <=  32'b00000000000000000000000000000000 ;
        335:  q   <=  32'b00000000000000000000000000000000 ;
        336:  q   <=  32'b00000000000000000000000000000000 ;
        337:  q   <=  32'b00000000000000000000000000000000 ;
        338:  q   <=  32'b00000000000000000000000000000000 ;
        339:  q   <=  32'b00000000000000000000000000000000 ;
        340:  q   <=  32'b00000000000000000000000000000000 ;
        341:  q   <=  32'b00000000000000000000000000000000 ;
        342:  q   <=  32'b00000000000000000000000000000000 ;
        343:  q   <=  32'b00000000000000000000000000000000 ;
        344:  q   <=  32'b00000000000000000000000000000000 ;
        345:  q   <=  32'b00000000000000000000000000000000 ;
        346:  q   <=  32'b00000000000000000000000000000000 ;
        347:  q   <=  32'b00000000000000000000000000000000 ;
        348:  q   <=  32'b00000000000000000000000000000000 ;
        349:  q   <=  32'b00000000000000000000000000000000 ;
        350:  q   <=  32'b00000000000000000000000000000000 ;
        351:  q   <=  32'b00000000000000000000000000000000 ;
        352:  q   <=  32'b00000000000000000000000000000000 ;
        353:  q   <=  32'b00000000000000000000000000000000 ;
        354:  q   <=  32'b00000000000000000000000000000000 ;
        355:  q   <=  32'b00000000000000000000000000000000 ;
        356:  q   <=  32'b00000000000000000000000000000000 ;
        357:  q   <=  32'b00000000000000000000000000000000 ;
        358:  q   <=  32'b00000000000000000000000000000000 ;
        359:  q   <=  32'b00000000000000000000000000000000 ;
        360:  q   <=  32'b00000000000000000000000000000000 ;
        361:  q   <=  32'b00000000000000000000000000000000 ;
        362:  q   <=  32'b00000000000000000000000000000000 ;
        363:  q   <=  32'b00000000000000000000000000000000 ;
        364:  q   <=  32'b00000000000000000000000000000000 ;
        365:  q   <=  32'b00000000000000000000000000000000 ;
        366:  q   <=  32'b00000000000000000000000000000000 ;
        367:  q   <=  32'b00000000000000000000000000000000 ;
        368:  q   <=  32'b00000000000000000000000000000000 ;
        369:  q   <=  32'b00000000000000000000000000000000 ;
        370:  q   <=  32'b00000000000000000000000000000000 ;
        371:  q   <=  32'b00000000000000000000000000000000 ;
        372:  q   <=  32'b00000000000000000000000000000000 ;
        373:  q   <=  32'b00000000000000000000000000000000 ;
        374:  q   <=  32'b00000000000000000000000000000000 ;
        375:  q   <=  32'b00000000000000000000000000000000 ;
        376:  q   <=  32'b00000000000000000000000000000000 ;
        377:  q   <=  32'b00000000000000000000000000000000 ;
        378:  q   <=  32'b00000000000000000000000000000000 ;
        379:  q   <=  32'b00000000000000000000000000000000 ;
        380:  q   <=  32'b00000000000000000000000000000000 ;
        381:  q   <=  32'b00000000000000000000000000000000 ;
        382:  q   <=  32'b00000000000000000000000000000000 ;
        383:  q   <=  32'b00000000000000000000000000000000 ;
        384:  q   <=  32'b00000000000000000000000000000000 ;
        385:  q   <=  32'b00000000000000000000000000000000 ;
        386:  q   <=  32'b00000000000000000000000000000000 ;
        387:  q   <=  32'b00000000000000000000000000000000 ;
        388:  q   <=  32'b00000000000000000000000000000000 ;
        389:  q   <=  32'b00000000000000000000000000000000 ;
        390:  q   <=  32'b00000000000000000000000000000000 ;
        391:  q   <=  32'b00000000000000000000000000000000 ;
        392:  q   <=  32'b00111110101011010001010000110011 ;
        393:  q   <=  32'b00111111001100101000001011100001 ;
        394:  q   <=  32'b00111111100001101110010001110101 ;
        395:  q   <=  32'b00111111101101000010111100011101 ;
        396:  q   <=  32'b00111111111000010010001001101000 ;
        397:  q   <=  32'b00111111111100100100000010101101 ;
        398:  q   <=  32'b00111111110001011111100100101011 ;
        399:  q   <=  32'b00111111100110100000011000011110 ;
        400:  q   <=  32'b00111111010111001100110100101000 ;
        401:  q   <=  32'b00111111000001100011001101000010 ;
        402:  q   <=  32'b00111110010000001111001011010110 ;
        403:  q   <=  32'b00000000000000000000000000000000 ;
        404:  q   <=  32'b00000000000000000000000000000000 ;
        405:  q   <=  32'b00000000000000000000000000000000 ;
        406:  q   <=  32'b00000000000000000000000000000000 ;
        407:  q   <=  32'b00000000000000000000000000000000 ;
        408:  q   <=  32'b00000000000000000000000000000000 ;
        409:  q   <=  32'b00000000000000000000000000000000 ;
        410:  q   <=  32'b00000000000000000000000000000000 ;
        411:  q   <=  32'b00000000000000000000000000000000 ;
        412:  q   <=  32'b00000000000000000000000000000000 ;
        413:  q   <=  32'b00000000000000000000000000000000 ;
        414:  q   <=  32'b00000000000000000000000000000000 ;
        415:  q   <=  32'b00000000000000000000000000000000 ;
        416:  q   <=  32'b00000000000000000000000000000000 ;
        417:  q   <=  32'b00000000000000000000000000000000 ;
        418:  q   <=  32'b00000000000000000000000000000000 ;
        419:  q   <=  32'b00000000000000000000000000000000 ;
        420:  q   <=  32'b00000000000000000000000000000000 ;
        421:  q   <=  32'b00000000000000000000000000000000 ;
        422:  q   <=  32'b00000000000000000000000000000000 ;
        423:  q   <=  32'b00000000000000000000000000000000 ;
        424:  q   <=  32'b00000000000000000000000000000000 ;
        425:  q   <=  32'b00000000000000000000000000000000 ;
        426:  q   <=  32'b00000000000000000000000000000000 ;
        427:  q   <=  32'b00000000000000000000000000000000 ;
        428:  q   <=  32'b00000000000000000000000000000000 ;
        429:  q   <=  32'b00000000000000000000000000000000 ;
        430:  q   <=  32'b00000000000000000000000000000000 ;
        431:  q   <=  32'b00000000000000000000000000000000 ;
        432:  q   <=  32'b00000000000000000000000000000000 ;
        433:  q   <=  32'b00000000000000000000000000000000 ;
        434:  q   <=  32'b00000000000000000000000000000000 ;
        435:  q   <=  32'b00000000000000000000000000000000 ;
        436:  q   <=  32'b00000000000000000000000000000000 ;
        437:  q   <=  32'b00000000000000000000000000000000 ;
        438:  q   <=  32'b00000000000000000000000000000000 ;
        439:  q   <=  32'b00000000000000000000000000000000 ;
        440:  q   <=  32'b00000000000000000000000000000000 ;
        441:  q   <=  32'b00000000000000000000000000000000 ;
        442:  q   <=  32'b00000000000000000000000000000000 ;
        443:  q   <=  32'b00000000000000000000000000000000 ;
        444:  q   <=  32'b00000000000000000000000000000000 ;
        445:  q   <=  32'b00000000000000000000000000000000 ;
        446:  q   <=  32'b00000000000000000000000000000000 ;
        447:  q   <=  32'b00000000000000000000000000000000 ;
        448:  q   <=  32'b00000000000000000000000000000000 ;
        449:  q   <=  32'b00000000000000000000000000000000 ;
        450:  q   <=  32'b00000000000000000000000000000000 ;
        451:  q   <=  32'b00000000000000000000000000000000 ;
        452:  q   <=  32'b00000000000000000000000000000000 ;
        453:  q   <=  32'b00000000000000000000000000000000 ;
        454:  q   <=  32'b00000000000000000000000000000000 ;
        455:  q   <=  32'b00000000000000000000000000000000 ;
        456:  q   <=  32'b00000000000000000000000000000000 ;
        457:  q   <=  32'b00000000000000000000000000000000 ;
        458:  q   <=  32'b00000000000000000000000000000000 ;
        459:  q   <=  32'b00000000000000000000000000000000 ;
        460:  q   <=  32'b00000000000000000000000000000000 ;
        461:  q   <=  32'b00000000000000000000000000000000 ;
        462:  q   <=  32'b00000000000000000000000000000000 ;
        463:  q   <=  32'b00000000000000000000000000000000 ;
        464:  q   <=  32'b00000000000000000000000000000000 ;
        465:  q   <=  32'b00000000000000000000000000000000 ;
        466:  q   <=  32'b00000000000000000000000000000000 ;
        467:  q   <=  32'b00000000000000000000000000000000 ;
        468:  q   <=  32'b00000000000000000000000000000000 ;
        469:  q   <=  32'b00000000000000000000000000000000 ;
        470:  q   <=  32'b00000000000000000000000000000000 ;
        471:  q   <=  32'b00000000000000000000000000000000 ;
        472:  q   <=  32'b00000000000000000000000000000000 ;
        473:  q   <=  32'b00000000000000000000000000000000 ;
        474:  q   <=  32'b00000000000000000000000000000000 ;
        475:  q   <=  32'b00000000000000000000000000000000 ;
        476:  q   <=  32'b00000000000000000000000000000000 ;
        477:  q   <=  32'b00000000000000000000000000000000 ;
        478:  q   <=  32'b00000000000000000000000000000000 ;
        479:  q   <=  32'b00000000000000000000000000000000 ;
        480:  q   <=  32'b00000000000000000000000000000000 ;
        481:  q   <=  32'b00000000000000000000000000000000 ;
        482:  q   <=  32'b00000000000000000000000000000000 ;
        483:  q   <=  32'b00000000000000000000000000000000 ;
        484:  q   <=  32'b00000000000000000000000000000000 ;
        485:  q   <=  32'b00000000000000000000000000000000 ;
        486:  q   <=  32'b00000000000000000000000000000000 ;
        487:  q   <=  32'b00000000000000000000000000000000 ;
        488:  q   <=  32'b00000000000000000000000000000000 ;
        489:  q   <=  32'b00000000000000000000000000000000 ;
        490:  q   <=  32'b00000000000000000000000000000000 ;
        491:  q   <=  32'b00000000000000000000000000000000 ;
        492:  q   <=  32'b00000000000000000000000000000000 ;
        493:  q   <=  32'b00000000000000000000000000000000 ;
        494:  q   <=  32'b00000000000000000000000000000000 ;
        495:  q   <=  32'b00000000000000000000000000000000 ;
        496:  q   <=  32'b00000000000000000000000000000000 ;
        497:  q   <=  32'b00000000000000000000000000000000 ;
        498:  q   <=  32'b00000000000000000000000000000000 ;
        499:  q   <=  32'b00000000000000000000000000000000 ;
        500:  q   <=  32'b00000000000000000000000000000000 ;
        501:  q   <=  32'b00000000000000000000000000000000 ;
        502:  q   <=  32'b00000000000000000000000000000000 ;
        503:  q   <=  32'b00000000000000000000000000000000 ;
        504:  q   <=  32'b00000000000000000000000000000000 ;
        505:  q   <=  32'b00000000000000000000000000000000 ;
        506:  q   <=  32'b00000000000000000000000000000000 ;
        507:  q   <=  32'b00000000000000000000000000000000 ;
        508:  q   <=  32'b00000000000000000000000000000000 ;
        509:  q   <=  32'b00000000000000000000000000000000 ;
        510:  q   <=  32'b00000000000000000000000000000000 ;
        511:  q   <=  32'b00000000000000000000000000000000 ;
        512:  q   <=  32'b00000000000000000000000000000000 ;
        513:  q   <=  32'b00000000000000000000000000000000 ;
        514:  q   <=  32'b00000000000000000000000000000000 ;
        515:  q   <=  32'b00000000000000000000000000000000 ;
        516:  q   <=  32'b00000000000000000000000000000000 ;
        517:  q   <=  32'b00000000000000000000000000000000 ;
        518:  q   <=  32'b00000000000000000000000000000000 ;
        519:  q   <=  32'b00000000000000000000000000000000 ;
        520:  q   <=  32'b00000000000000000000000000000000 ;
        521:  q   <=  32'b00000000000000000000000000000000 ;
        522:  q   <=  32'b00000000000000000000000000000000 ;
        523:  q   <=  32'b00000000000000000000000000000000 ;
        524:  q   <=  32'b00000000000000000000000000000000 ;
        525:  q   <=  32'b00000000000000000000000000000000 ;
        526:  q   <=  32'b00000000000000000000000000000000 ;
        527:  q   <=  32'b00000000000000000000000000000000 ;
        528:  q   <=  32'b00000000000000000000000000000000 ;
        529:  q   <=  32'b00000000000000000000000000000000 ;
        530:  q   <=  32'b00000000000000000000000000000000 ;
        531:  q   <=  32'b00000000000000000000000000000000 ;
        532:  q   <=  32'b00000000000000000000000000000000 ;
        533:  q   <=  32'b00000000000000000000000000000000 ;
        534:  q   <=  32'b00000000000000000000000000000000 ;
        535:  q   <=  32'b00000000000000000000000000000000 ;
        536:  q   <=  32'b00000000000000000000000000000000 ;
        537:  q   <=  32'b00000000000000000000000000000000 ;
        538:  q   <=  32'b00000000000000000000000000000000 ;
        539:  q   <=  32'b00000000000000000000000000000000 ;
        540:  q   <=  32'b00000000000000000000000000000000 ;
        541:  q   <=  32'b00000000000000000000000000000000 ;
        542:  q   <=  32'b00000000000000000000000000000000 ;
        543:  q   <=  32'b00000000000000000000000000000000 ;
        544:  q   <=  32'b00000000000000000000000000000000 ;
        545:  q   <=  32'b00000000000000000000000000000000 ;
        546:  q   <=  32'b00000000000000000000000000000000 ;
        547:  q   <=  32'b00000000000000000000000000000000 ;
        548:  q   <=  32'b00000000000000000000000000000000 ;
        549:  q   <=  32'b00000000000000000000000000000000 ;
        550:  q   <=  32'b00000000000000000000000000000000 ;
        551:  q   <=  32'b00000000000000000000000000000000 ;
        552:  q   <=  32'b00000000000000000000000000000000 ;
        553:  q   <=  32'b00000000000000000000000000000000 ;
        554:  q   <=  32'b00000000000000000000000000000000 ;
        555:  q   <=  32'b00000000000000000000000000000000 ;
        556:  q   <=  32'b00000000000000000000000000000000 ;
        557:  q   <=  32'b00000000000000000000000000000000 ;
        558:  q   <=  32'b00000000000000000000000000000000 ;
        559:  q   <=  32'b00000000000000000000000000000000 ;
        560:  q   <=  32'b00000000000000000000000000000000 ;
        561:  q   <=  32'b00000000000000000000000000000000 ;
        562:  q   <=  32'b00000000000000000000000000000000 ;
        563:  q   <=  32'b00000000000000000000000000000000 ;
        564:  q   <=  32'b00000000000000000000000000000000 ;
        565:  q   <=  32'b00000000000000000000000000000000 ;
        566:  q   <=  32'b00000000000000000000000000000000 ;
        567:  q   <=  32'b00000000000000000000000000000000 ;
        568:  q   <=  32'b00000000000000000000000000000000 ;
        569:  q   <=  32'b00000000000000000000000000000000 ;
        570:  q   <=  32'b00000000000000000000000000000000 ;
        571:  q   <=  32'b00000000000000000000000000000000 ;
        572:  q   <=  32'b00000000000000000000000000000000 ;
        573:  q   <=  32'b00000000000000000000000000000000 ;
        574:  q   <=  32'b00000000000000000000000000000000 ;
        575:  q   <=  32'b00000000000000000000000000000000 ;
        576:  q   <=  32'b00000000000000000000000000000000 ;
        577:  q   <=  32'b00000000000000000000000000000000 ;
        578:  q   <=  32'b00000000000000000000000000000000 ;
        579:  q   <=  32'b00000000000000000000000000000000 ;
        580:  q   <=  32'b00000000000000000000000000000000 ;
        581:  q   <=  32'b00000000000000000000000000000000 ;
        582:  q   <=  32'b00000000000000000000000000000000 ;
        583:  q   <=  32'b00000000000000000000000000000000 ;
        584:  q   <=  32'b00000000000000000000000000000000 ;
        585:  q   <=  32'b00000000000000000000000000000000 ;
        586:  q   <=  32'b00000000000000000000000000000000 ;
        587:  q   <=  32'b00000000000000000000000000000000 ;
        588:  q   <=  32'b00000000000000000000000000000000 ;
        589:  q   <=  32'b00000000000000000000000000000000 ;
        590:  q   <=  32'b00000000000000000000000000000000 ;
        591:  q   <=  32'b00000000000000000000000000000000 ;
        592:  q   <=  32'b00000000000000000000000000000000 ;
        593:  q   <=  32'b00000000000000000000000000000000 ;
        594:  q   <=  32'b00000000000000000000000000000000 ;
        595:  q   <=  32'b00000000000000000000000000000000 ;
        596:  q   <=  32'b00000000000000000000000000000000 ;
        597:  q   <=  32'b00000000000000000000000000000000 ;
        598:  q   <=  32'b00000000000000000000000000000000 ;
        599:  q   <=  32'b00000000000000000000000000000000 ;
        600:  q   <=  32'b00000000000000000000000000000000 ;
        601:  q   <=  32'b00000000000000000000000000000000 ;
        602:  q   <=  32'b00000000000000000000000000000000 ;
        603:  q   <=  32'b00000000000000000000000000000000 ;
        604:  q   <=  32'b00000000000000000000000000000000 ;
        605:  q   <=  32'b00000000000000000000000000000000 ;
        606:  q   <=  32'b00000000000000000000000000000000 ;
        607:  q   <=  32'b00000000000000000000000000000000 ;
        608:  q   <=  32'b00000000000000000000000000000000 ;
        609:  q   <=  32'b00000000000000000000000000000000 ;
        610:  q   <=  32'b00000000000000000000000000000000 ;
        611:  q   <=  32'b00000000000000000000000000000000 ;
        612:  q   <=  32'b00000000000000000000000000000000 ;
        613:  q   <=  32'b00000000000000000000000000000000 ;
        614:  q   <=  32'b00000000000000000000000000000000 ;
        615:  q   <=  32'b00000000000000000000000000000000 ;
        616:  q   <=  32'b00000000000000000000000000000000 ;
        617:  q   <=  32'b00000000000000000000000000000000 ;
        618:  q   <=  32'b00000000000000000000000000000000 ;
        619:  q   <=  32'b00000000000000000000000000000000 ;
        620:  q   <=  32'b00000000000000000000000000000000 ;
        621:  q   <=  32'b00000000000000000000000000000000 ;
        622:  q   <=  32'b00000000000000000000000000000000 ;
        623:  q   <=  32'b00000000000000000000000000000000 ;
        624:  q   <=  32'b00000000000000000000000000000000 ;
        625:  q   <=  32'b00000000000000000000000000000000 ;
        626:  q   <=  32'b00000000000000000000000000000000 ;
        627:  q   <=  32'b00000000000000000000000000000000 ;
        628:  q   <=  32'b00000000000000000000000000000000 ;
        629:  q   <=  32'b00000000000000000000000000000000 ;
        630:  q   <=  32'b00000000000000000000000000000000 ;
        631:  q   <=  32'b00000000000000000000000000000000 ;
        632:  q   <=  32'b00000000000000000000000000000000 ;
        633:  q   <=  32'b00000000000000000000000000000000 ;
        634:  q   <=  32'b00000000000000000000000000000000 ;
        635:  q   <=  32'b00000000000000000000000000000000 ;
        636:  q   <=  32'b00000000000000000000000000000000 ;
        637:  q   <=  32'b00000000000000000000000000000000 ;
        638:  q   <=  32'b00000000000000000000000000000000 ;
        639:  q   <=  32'b00000000000000000000000000000000 ;
        640:  q   <=  32'b00000000000000000000000000000000 ;
        641:  q   <=  32'b00000000000000000000000000000000 ;
        642:  q   <=  32'b00000000000000000000000000000000 ;
        643:  q   <=  32'b00000000000000000000000000000000 ;
        644:  q   <=  32'b00000000000000000000000000000000 ;
        645:  q   <=  32'b00000000000000000000000000000000 ;
        646:  q   <=  32'b00000000000000000000000000000000 ;
        647:  q   <=  32'b00000000000000000000000000000000 ;
        648:  q   <=  32'b00000000000000000000000000000000 ;
        649:  q   <=  32'b00000000000000000000000000000000 ;
        650:  q   <=  32'b00000000000000000000000000000000 ;
        651:  q   <=  32'b00000000000000000000000000000000 ;
        652:  q   <=  32'b00000000000000000000000000000000 ;
        653:  q   <=  32'b00111101110110111111010100101101 ;
        654:  q   <=  32'b00111110111010000001101101010010 ;
        655:  q   <=  32'b00111111010010111111001111000011 ;
        656:  q   <=  32'b00111111100100011001100101101011 ;
        657:  q   <=  32'b00111111101111001110011001011110 ;
        658:  q   <=  32'b00111111111001111110000110100101 ;
        659:  q   <=  32'b00111111111011010111001111011011 ;
        660:  q   <=  32'b00111111110000110001100100111111 ;
        661:  q   <=  32'b00111111100110010000110110100111 ;
        662:  q   <=  32'b00111111010111101010000001101110 ;
        663:  q   <=  32'b00111111000010111100000000101011 ;
        664:  q   <=  32'b00111110011001011110001101101001 ;
        665:  q   <=  32'b00000000000000000000000000000000 ;
        666:  q   <=  32'b00000000000000000000000000000000 ;
        667:  q   <=  32'b00000000000000000000000000000000 ;
        668:  q   <=  32'b00000000000000000000000000000000 ;
        669:  q   <=  32'b00000000000000000000000000000000 ;
        670:  q   <=  32'b00000000000000000000000000000000 ;
        671:  q   <=  32'b00000000000000000000000000000000 ;
        672:  q   <=  32'b00000000000000000000000000000000 ;
        673:  q   <=  32'b00000000000000000000000000000000 ;
        674:  q   <=  32'b00000000000000000000000000000000 ;
        675:  q   <=  32'b00000000000000000000000000000000 ;
        676:  q   <=  32'b00000000000000000000000000000000 ;
        677:  q   <=  32'b00000000000000000000000000000000 ;
        678:  q   <=  32'b00000000000000000000000000000000 ;
        679:  q   <=  32'b00000000000000000000000000000000 ;
        680:  q   <=  32'b00000000000000000000000000000000 ;
        681:  q   <=  32'b00000000000000000000000000000000 ;
        682:  q   <=  32'b00000000000000000000000000000000 ;
        683:  q   <=  32'b00000000000000000000000000000000 ;
        684:  q   <=  32'b00000000000000000000000000000000 ;
        685:  q   <=  32'b00000000000000000000000000000000 ;
        686:  q   <=  32'b00000000000000000000000000000000 ;
        687:  q   <=  32'b00000000000000000000000000000000 ;
        688:  q   <=  32'b00000000000000000000000000000000 ;
        689:  q   <=  32'b00000000000000000000000000000000 ;
        690:  q   <=  32'b00000000000000000000000000000000 ;
        691:  q   <=  32'b00000000000000000000000000000000 ;
        692:  q   <=  32'b00000000000000000000000000000000 ;
        693:  q   <=  32'b00000000000000000000000000000000 ;
        694:  q   <=  32'b00000000000000000000000000000000 ;
        695:  q   <=  32'b00000000000000000000000000000000 ;
        696:  q   <=  32'b00000000000000000000000000000000 ;
        697:  q   <=  32'b00000000000000000000000000000000 ;
        698:  q   <=  32'b00000000000000000000000000000000 ;
        699:  q   <=  32'b00000000000000000000000000000000 ;
        700:  q   <=  32'b00000000000000000000000000000000 ;
        701:  q   <=  32'b00000000000000000000000000000000 ;
        702:  q   <=  32'b00000000000000000000000000000000 ;
        703:  q   <=  32'b00000000000000000000000000000000 ;
        704:  q   <=  32'b00000000000000000000000000000000 ;
        705:  q   <=  32'b00000000000000000000000000000000 ;
        706:  q   <=  32'b00000000000000000000000000000000 ;
        707:  q   <=  32'b00000000000000000000000000000000 ;
        708:  q   <=  32'b00000000000000000000000000000000 ;
        709:  q   <=  32'b00000000000000000000000000000000 ;
        710:  q   <=  32'b00000000000000000000000000000000 ;
        711:  q   <=  32'b00000000000000000000000000000000 ;
        712:  q   <=  32'b00000000000000000000000000000000 ;
        713:  q   <=  32'b00000000000000000000000000000000 ;
        714:  q   <=  32'b00000000000000000000000000000000 ;
        715:  q   <=  32'b00000000000000000000000000000000 ;
        716:  q   <=  32'b00000000000000000000000000000000 ;
        717:  q   <=  32'b00000000000000000000000000000000 ;
        718:  q   <=  32'b00000000000000000000000000000000 ;
        719:  q   <=  32'b00000000000000000000000000000000 ;
        720:  q   <=  32'b00000000000000000000000000000000 ;
        721:  q   <=  32'b00000000000000000000000000000000 ;
        722:  q   <=  32'b00000000000000000000000000000000 ;
        723:  q   <=  32'b00000000000000000000000000000000 ;
        724:  q   <=  32'b00000000000000000000000000000000 ;
        725:  q   <=  32'b00000000000000000000000000000000 ;
        726:  q   <=  32'b00000000000000000000000000000000 ;
        727:  q   <=  32'b00000000000000000000000000000000 ;
        728:  q   <=  32'b00000000000000000000000000000000 ;
        729:  q   <=  32'b00000000000000000000000000000000 ;
        730:  q   <=  32'b00000000000000000000000000000000 ;
        731:  q   <=  32'b00000000000000000000000000000000 ;
        732:  q   <=  32'b00000000000000000000000000000000 ;
        733:  q   <=  32'b00000000000000000000000000000000 ;
        734:  q   <=  32'b00000000000000000000000000000000 ;
        735:  q   <=  32'b00000000000000000000000000000000 ;
        736:  q   <=  32'b00000000000000000000000000000000 ;
        737:  q   <=  32'b00000000000000000000000000000000 ;
        738:  q   <=  32'b00000000000000000000000000000000 ;
        739:  q   <=  32'b00000000000000000000000000000000 ;
        740:  q   <=  32'b00000000000000000000000000000000 ;
        741:  q   <=  32'b00000000000000000000000000000000 ;
        742:  q   <=  32'b00000000000000000000000000000000 ;
        743:  q   <=  32'b00000000000000000000000000000000 ;
        744:  q   <=  32'b00000000000000000000000000000000 ;
        745:  q   <=  32'b00000000000000000000000000000000 ;
        746:  q   <=  32'b00000000000000000000000000000000 ;
        747:  q   <=  32'b00000000000000000000000000000000 ;
        748:  q   <=  32'b00000000000000000000000000000000 ;
        749:  q   <=  32'b00000000000000000000000000000000 ;
        750:  q   <=  32'b00000000000000000000000000000000 ;
        751:  q   <=  32'b00000000000000000000000000000000 ;
        752:  q   <=  32'b00000000000000000000000000000000 ;
        753:  q   <=  32'b00000000000000000000000000000000 ;
        754:  q   <=  32'b00000000000000000000000000000000 ;
        755:  q   <=  32'b00000000000000000000000000000000 ;
        756:  q   <=  32'b00000000000000000000000000000000 ;
        757:  q   <=  32'b00000000000000000000000000000000 ;
        758:  q   <=  32'b00000000000000000000000000000000 ;
        759:  q   <=  32'b00000000000000000000000000000000 ;
        760:  q   <=  32'b00000000000000000000000000000000 ;
        761:  q   <=  32'b00000000000000000000000000000000 ;
        762:  q   <=  32'b00000000000000000000000000000000 ;
        763:  q   <=  32'b00000000000000000000000000000000 ;
        764:  q   <=  32'b00000000000000000000000000000000 ;
        765:  q   <=  32'b00000000000000000000000000000000 ;
        766:  q   <=  32'b00000000000000000000000000000000 ;
        767:  q   <=  32'b00000000000000000000000000000000 ;
        768:  q   <=  32'b00000000000000000000000000000000 ;
        769:  q   <=  32'b00000000000000000000000000000000 ;
        770:  q   <=  32'b00000000000000000000000000000000 ;
        771:  q   <=  32'b00000000000000000000000000000000 ;
        772:  q   <=  32'b00000000000000000000000000000000 ;
        773:  q   <=  32'b00000000000000000000000000000000 ;
        774:  q   <=  32'b00000000000000000000000000000000 ;
        775:  q   <=  32'b00000000000000000000000000000000 ;
        776:  q   <=  32'b00000000000000000000000000000000 ;
        777:  q   <=  32'b00000000000000000000000000000000 ;
        778:  q   <=  32'b00000000000000000000000000000000 ;
        779:  q   <=  32'b00000000000000000000000000000000 ;
        780:  q   <=  32'b00000000000000000000000000000000 ;
        781:  q   <=  32'b00000000000000000000000000000000 ;
        782:  q   <=  32'b00000000000000000000000000000000 ;
        783:  q   <=  32'b00000000000000000000000000000000 ;
        784:  q   <=  32'b00000000000000000000000000000000 ;
        785:  q   <=  32'b00000000000000000000000000000000 ;
        786:  q   <=  32'b00000000000000000000000000000000 ;
        787:  q   <=  32'b00000000000000000000000000000000 ;
        788:  q   <=  32'b00000000000000000000000000000000 ;
        789:  q   <=  32'b00000000000000000000000000000000 ;
        790:  q   <=  32'b00000000000000000000000000000000 ;
        791:  q   <=  32'b00000000000000000000000000000000 ;
        792:  q   <=  32'b00000000000000000000000000000000 ;
        793:  q   <=  32'b00000000000000000000000000000000 ;
        794:  q   <=  32'b00000000000000000000000000000000 ;
        795:  q   <=  32'b00000000000000000000000000000000 ;
        796:  q   <=  32'b00000000000000000000000000000000 ;
        797:  q   <=  32'b00000000000000000000000000000000 ;
        798:  q   <=  32'b00000000000000000000000000000000 ;
        799:  q   <=  32'b00000000000000000000000000000000 ;
        800:  q   <=  32'b00000000000000000000000000000000 ;
        801:  q   <=  32'b00000000000000000000000000000000 ;
        802:  q   <=  32'b00000000000000000000000000000000 ;
        803:  q   <=  32'b00000000000000000000000000000000 ;
        804:  q   <=  32'b00000000000000000000000000000000 ;
        805:  q   <=  32'b00000000000000000000000000000000 ;
        806:  q   <=  32'b00000000000000000000000000000000 ;
        807:  q   <=  32'b00000000000000000000000000000000 ;
        808:  q   <=  32'b00000000000000000000000000000000 ;
        809:  q   <=  32'b00000000000000000000000000000000 ;
        810:  q   <=  32'b00000000000000000000000000000000 ;
        811:  q   <=  32'b00000000000000000000000000000000 ;
        812:  q   <=  32'b00000000000000000000000000000000 ;
        813:  q   <=  32'b00000000000000000000000000000000 ;
        814:  q   <=  32'b00000000000000000000000000000000 ;
        815:  q   <=  32'b00000000000000000000000000000000 ;
        816:  q   <=  32'b00000000000000000000000000000000 ;
        817:  q   <=  32'b00000000000000000000000000000000 ;
        818:  q   <=  32'b00000000000000000000000000000000 ;
        819:  q   <=  32'b00000000000000000000000000000000 ;
        820:  q   <=  32'b00000000000000000000000000000000 ;
        821:  q   <=  32'b00000000000000000000000000000000 ;
        822:  q   <=  32'b00000000000000000000000000000000 ;
        823:  q   <=  32'b00000000000000000000000000000000 ;
        824:  q   <=  32'b00000000000000000000000000000000 ;
        825:  q   <=  32'b00000000000000000000000000000000 ;
        826:  q   <=  32'b00000000000000000000000000000000 ;
        827:  q   <=  32'b00000000000000000000000000000000 ;
        828:  q   <=  32'b00000000000000000000000000000000 ;
        829:  q   <=  32'b00000000000000000000000000000000 ;
        830:  q   <=  32'b00000000000000000000000000000000 ;
        831:  q   <=  32'b00000000000000000000000000000000 ;
        832:  q   <=  32'b00000000000000000000000000000000 ;
        833:  q   <=  32'b00000000000000000000000000000000 ;
        834:  q   <=  32'b00000000000000000000000000000000 ;
        835:  q   <=  32'b00000000000000000000000000000000 ;
        836:  q   <=  32'b00000000000000000000000000000000 ;
        837:  q   <=  32'b00000000000000000000000000000000 ;
        838:  q   <=  32'b00000000000000000000000000000000 ;
        839:  q   <=  32'b00000000000000000000000000000000 ;
        840:  q   <=  32'b00000000000000000000000000000000 ;
        841:  q   <=  32'b00000000000000000000000000000000 ;
        842:  q   <=  32'b00000000000000000000000000000000 ;
        843:  q   <=  32'b00000000000000000000000000000000 ;
        844:  q   <=  32'b00000000000000000000000000000000 ;
        845:  q   <=  32'b00000000000000000000000000000000 ;
        846:  q   <=  32'b00000000000000000000000000000000 ;
        847:  q   <=  32'b00000000000000000000000000000000 ;
        848:  q   <=  32'b00000000000000000000000000000000 ;
        849:  q   <=  32'b00000000000000000000000000000000 ;
        850:  q   <=  32'b00000000000000000000000000000000 ;
        851:  q   <=  32'b00000000000000000000000000000000 ;
        852:  q   <=  32'b00000000000000000000000000000000 ;
        853:  q   <=  32'b00000000000000000000000000000000 ;
        854:  q   <=  32'b00000000000000000000000000000000 ;
        855:  q   <=  32'b00000000000000000000000000000000 ;
        856:  q   <=  32'b00000000000000000000000000000000 ;
        857:  q   <=  32'b00000000000000000000000000000000 ;
        858:  q   <=  32'b00000000000000000000000000000000 ;
        859:  q   <=  32'b00000000000000000000000000000000 ;
        860:  q   <=  32'b00000000000000000000000000000000 ;
        861:  q   <=  32'b00000000000000000000000000000000 ;
        862:  q   <=  32'b00000000000000000000000000000000 ;
        863:  q   <=  32'b00000000000000000000000000000000 ;
        864:  q   <=  32'b00000000000000000000000000000000 ;
        865:  q   <=  32'b00000000000000000000000000000000 ;
        866:  q   <=  32'b00000000000000000000000000000000 ;
        867:  q   <=  32'b00000000000000000000000000000000 ;
        868:  q   <=  32'b00000000000000000000000000000000 ;
        869:  q   <=  32'b00000000000000000000000000000000 ;
        870:  q   <=  32'b00000000000000000000000000000000 ;
        871:  q   <=  32'b00000000000000000000000000000000 ;
        872:  q   <=  32'b00000000000000000000000000000000 ;
        873:  q   <=  32'b00000000000000000000000000000000 ;
        874:  q   <=  32'b00000000000000000000000000000000 ;
        875:  q   <=  32'b00000000000000000000000000000000 ;
        876:  q   <=  32'b00000000000000000000000000000000 ;
        877:  q   <=  32'b00000000000000000000000000000000 ;
        878:  q   <=  32'b00000000000000000000000000000000 ;
        879:  q   <=  32'b00000000000000000000000000000000 ;
        880:  q   <=  32'b00000000000000000000000000000000 ;
        881:  q   <=  32'b00000000000000000000000000000000 ;
        882:  q   <=  32'b00000000000000000000000000000000 ;
        883:  q   <=  32'b00000000000000000000000000000000 ;
        884:  q   <=  32'b00000000000000000000000000000000 ;
        885:  q   <=  32'b00000000000000000000000000000000 ;
        886:  q   <=  32'b00000000000000000000000000000000 ;
        887:  q   <=  32'b00000000000000000000000000000000 ;
        888:  q   <=  32'b00000000000000000000000000000000 ;
        889:  q   <=  32'b00000000000000000000000000000000 ;
        890:  q   <=  32'b00000000000000000000000000000000 ;
        891:  q   <=  32'b00000000000000000000000000000000 ;
        892:  q   <=  32'b00000000000000000000000000000000 ;
        893:  q   <=  32'b00000000000000000000000000000000 ;
        894:  q   <=  32'b00000000000000000000000000000000 ;
        895:  q   <=  32'b00000000000000000000000000000000 ;
        896:  q   <=  32'b00000000000000000000000000000000 ;
        897:  q   <=  32'b00000000000000000000000000000000 ;
        898:  q   <=  32'b00000000000000000000000000000000 ;
        899:  q   <=  32'b00000000000000000000000000000000 ;
        900:  q   <=  32'b00000000000000000000000000000000 ;
        901:  q   <=  32'b00000000000000000000000000000000 ;
        902:  q   <=  32'b00000000000000000000000000000000 ;
        903:  q   <=  32'b00000000000000000000000000000000 ;
        904:  q   <=  32'b00000000000000000000000000000000 ;
        905:  q   <=  32'b00000000000000000000000000000000 ;
        906:  q   <=  32'b00000000000000000000000000000000 ;
        907:  q   <=  32'b00000000000000000000000000000000 ;
        908:  q   <=  32'b00000000000000000000000000000000 ;
        909:  q   <=  32'b00000000000000000000000000000000 ;
        910:  q   <=  32'b00000000000000000000000000000000 ;
        911:  q   <=  32'b00000000000000000000000000000000 ;
        912:  q   <=  32'b00000000000000000000000000000000 ;
        913:  q   <=  32'b00000000000000000000000000000000 ;
        914:  q   <=  32'b00000000000000000000000000000000 ;
        915:  q   <=  32'b00111110000101000110000100100111 ;
        916:  q   <=  32'b00111110111100111001101100000011 ;
        917:  q   <=  32'b00111111010011011110010010110001 ;
        918:  q   <=  32'b00111111100100001010111111001000 ;
        919:  q   <=  32'b00111111101110100001111111101010 ;
        920:  q   <=  32'b00111111111000110100001110010010 ;
        921:  q   <=  32'b00111111111100111110010001101010 ;
        922:  q   <=  32'b00111111110010110101011100111101 ;
        923:  q   <=  32'b00111111101000110001010000011001 ;
        924:  q   <=  32'b00111111011101100011010001101000 ;
        925:  q   <=  32'b00111111001001101101000110001110 ;
        926:  q   <=  32'b00111110101011111111110000110100 ;
        927:  q   <=  32'b00111101000110111000100010011100 ;
        928:  q   <=  32'b00000000000000000000000000000000 ;
        929:  q   <=  32'b00000000000000000000000000000000 ;
        930:  q   <=  32'b00000000000000000000000000000000 ;
        931:  q   <=  32'b00000000000000000000000000000000 ;
        932:  q   <=  32'b00000000000000000000000000000000 ;
        933:  q   <=  32'b00000000000000000000000000000000 ;
        934:  q   <=  32'b00000000000000000000000000000000 ;
        935:  q   <=  32'b00000000000000000000000000000000 ;
        936:  q   <=  32'b00000000000000000000000000000000 ;
        937:  q   <=  32'b00000000000000000000000000000000 ;
        938:  q   <=  32'b00000000000000000000000000000000 ;
        939:  q   <=  32'b00000000000000000000000000000000 ;
        940:  q   <=  32'b00000000000000000000000000000000 ;
        941:  q   <=  32'b00000000000000000000000000000000 ;
        942:  q   <=  32'b00000000000000000000000000000000 ;
        943:  q   <=  32'b00000000000000000000000000000000 ;
        944:  q   <=  32'b00000000000000000000000000000000 ;
        945:  q   <=  32'b00000000000000000000000000000000 ;
        946:  q   <=  32'b00000000000000000000000000000000 ;
        947:  q   <=  32'b00000000000000000000000000000000 ;
        948:  q   <=  32'b00000000000000000000000000000000 ;
        949:  q   <=  32'b00000000000000000000000000000000 ;
        950:  q   <=  32'b00000000000000000000000000000000 ;
        951:  q   <=  32'b00000000000000000000000000000000 ;
        952:  q   <=  32'b00000000000000000000000000000000 ;
        953:  q   <=  32'b00000000000000000000000000000000 ;
        954:  q   <=  32'b00000000000000000000000000000000 ;
        955:  q   <=  32'b00000000000000000000000000000000 ;
        956:  q   <=  32'b00000000000000000000000000000000 ;
        957:  q   <=  32'b00000000000000000000000000000000 ;
        958:  q   <=  32'b00000000000000000000000000000000 ;
        959:  q   <=  32'b00000000000000000000000000000000 ;
        960:  q   <=  32'b00000000000000000000000000000000 ;
        961:  q   <=  32'b00000000000000000000000000000000 ;
        962:  q   <=  32'b00000000000000000000000000000000 ;
        963:  q   <=  32'b00000000000000000000000000000000 ;
        964:  q   <=  32'b00000000000000000000000000000000 ;
        965:  q   <=  32'b00000000000000000000000000000000 ;
        966:  q   <=  32'b00000000000000000000000000000000 ;
        967:  q   <=  32'b00000000000000000000000000000000 ;
        968:  q   <=  32'b00000000000000000000000000000000 ;
        969:  q   <=  32'b00000000000000000000000000000000 ;
        970:  q   <=  32'b00000000000000000000000000000000 ;
        971:  q   <=  32'b00000000000000000000000000000000 ;
        972:  q   <=  32'b00000000000000000000000000000000 ;
        973:  q   <=  32'b00000000000000000000000000000000 ;
        974:  q   <=  32'b00000000000000000000000000000000 ;
        975:  q   <=  32'b00000000000000000000000000000000 ;
        976:  q   <=  32'b00000000000000000000000000000000 ;
        977:  q   <=  32'b00000000000000000000000000000000 ;
        978:  q   <=  32'b00000000000000000000000000000000 ;
        979:  q   <=  32'b00000000000000000000000000000000 ;
        980:  q   <=  32'b00000000000000000000000000000000 ;
        981:  q   <=  32'b00000000000000000000000000000000 ;
        982:  q   <=  32'b00000000000000000000000000000000 ;
        983:  q   <=  32'b00000000000000000000000000000000 ;
        984:  q   <=  32'b00000000000000000000000000000000 ;
        985:  q   <=  32'b00000000000000000000000000000000 ;
        986:  q   <=  32'b00000000000000000000000000000000 ;
        987:  q   <=  32'b00000000000000000000000000000000 ;
        988:  q   <=  32'b00000000000000000000000000000000 ;
        989:  q   <=  32'b00000000000000000000000000000000 ;
        990:  q   <=  32'b00000000000000000000000000000000 ;
        991:  q   <=  32'b00000000000000000000000000000000 ;
        992:  q   <=  32'b00000000000000000000000000000000 ;
        993:  q   <=  32'b00000000000000000000000000000000 ;
        994:  q   <=  32'b00000000000000000000000000000000 ;
        995:  q   <=  32'b00000000000000000000000000000000 ;
        996:  q   <=  32'b00000000000000000000000000000000 ;
        997:  q   <=  32'b00000000000000000000000000000000 ;
        998:  q   <=  32'b00000000000000000000000000000000 ;
        999:  q   <=  32'b00000000000000000000000000000000 ;
        1000:  q   <=  32'b00000000000000000000000000000000 ;
        1001:  q   <=  32'b00000000000000000000000000000000 ;
        1002:  q   <=  32'b00000000000000000000000000000000 ;
        1003:  q   <=  32'b00000000000000000000000000000000 ;
        1004:  q   <=  32'b00000000000000000000000000000000 ;
        1005:  q   <=  32'b00000000000000000000000000000000 ;
        1006:  q   <=  32'b00000000000000000000000000000000 ;
        1007:  q   <=  32'b00000000000000000000000000000000 ;
        1008:  q   <=  32'b00000000000000000000000000000000 ;
        1009:  q   <=  32'b00000000000000000000000000000000 ;
        1010:  q   <=  32'b00000000000000000000000000000000 ;
        1011:  q   <=  32'b00000000000000000000000000000000 ;
        1012:  q   <=  32'b00000000000000000000000000000000 ;
        1013:  q   <=  32'b00000000000000000000000000000000 ;
        1014:  q   <=  32'b00000000000000000000000000000000 ;
        1015:  q   <=  32'b00000000000000000000000000000000 ;
        1016:  q   <=  32'b00000000000000000000000000000000 ;
        1017:  q   <=  32'b00000000000000000000000000000000 ;
        1018:  q   <=  32'b00000000000000000000000000000000 ;
        1019:  q   <=  32'b00000000000000000000000000000000 ;
        1020:  q   <=  32'b00000000000000000000000000000000 ;
        1021:  q   <=  32'b00000000000000000000000000000000 ;
        1022:  q   <=  32'b00000000000000000000000000000000 ;
        1023:  q   <=  32'b00000000000000000000000000000000 ;
        1024:  q   <=  32'b00000000000000000000000000000000 ;
        1025:  q   <=  32'b00000000000000000000000000000000 ;
        1026:  q   <=  32'b00000000000000000000000000000000 ;
        1027:  q   <=  32'b00000000000000000000000000000000 ;
        1028:  q   <=  32'b00000000000000000000000000000000 ;
        1029:  q   <=  32'b00000000000000000000000000000000 ;
        1030:  q   <=  32'b00000000000000000000000000000000 ;
        1031:  q   <=  32'b00000000000000000000000000000000 ;
        1032:  q   <=  32'b00000000000000000000000000000000 ;
        1033:  q   <=  32'b00000000000000000000000000000000 ;
        1034:  q   <=  32'b00000000000000000000000000000000 ;
        1035:  q   <=  32'b00000000000000000000000000000000 ;
        1036:  q   <=  32'b00000000000000000000000000000000 ;
        1037:  q   <=  32'b00000000000000000000000000000000 ;
        1038:  q   <=  32'b00000000000000000000000000000000 ;
        1039:  q   <=  32'b00000000000000000000000000000000 ;
        1040:  q   <=  32'b00000000000000000000000000000000 ;
        1041:  q   <=  32'b00000000000000000000000000000000 ;
        1042:  q   <=  32'b00000000000000000000000000000000 ;
        1043:  q   <=  32'b00000000000000000000000000000000 ;
        1044:  q   <=  32'b00000000000000000000000000000000 ;
        1045:  q   <=  32'b00000000000000000000000000000000 ;
        1046:  q   <=  32'b00000000000000000000000000000000 ;
        1047:  q   <=  32'b00000000000000000000000000000000 ;
        1048:  q   <=  32'b00000000000000000000000000000000 ;
        1049:  q   <=  32'b00000000000000000000000000000000 ;
        1050:  q   <=  32'b00000000000000000000000000000000 ;
        1051:  q   <=  32'b00000000000000000000000000000000 ;
        1052:  q   <=  32'b00000000000000000000000000000000 ;
        1053:  q   <=  32'b00000000000000000000000000000000 ;
        1054:  q   <=  32'b00000000000000000000000000000000 ;
        1055:  q   <=  32'b00000000000000000000000000000000 ;
        1056:  q   <=  32'b00000000000000000000000000000000 ;
        1057:  q   <=  32'b00000000000000000000000000000000 ;
        1058:  q   <=  32'b00000000000000000000000000000000 ;
        1059:  q   <=  32'b00000000000000000000000000000000 ;
        1060:  q   <=  32'b00000000000000000000000000000000 ;
        1061:  q   <=  32'b00000000000000000000000000000000 ;
        1062:  q   <=  32'b00000000000000000000000000000000 ;
        1063:  q   <=  32'b00000000000000000000000000000000 ;
        1064:  q   <=  32'b00000000000000000000000000000000 ;
        1065:  q   <=  32'b00000000000000000000000000000000 ;
        1066:  q   <=  32'b00000000000000000000000000000000 ;
        1067:  q   <=  32'b00000000000000000000000000000000 ;
        1068:  q   <=  32'b00000000000000000000000000000000 ;
        1069:  q   <=  32'b00000000000000000000000000000000 ;
        1070:  q   <=  32'b00000000000000000000000000000000 ;
        1071:  q   <=  32'b00000000000000000000000000000000 ;
        1072:  q   <=  32'b00000000000000000000000000000000 ;
        1073:  q   <=  32'b00000000000000000000000000000000 ;
        1074:  q   <=  32'b00000000000000000000000000000000 ;
        1075:  q   <=  32'b00000000000000000000000000000000 ;
        1076:  q   <=  32'b00000000000000000000000000000000 ;
        1077:  q   <=  32'b00000000000000000000000000000000 ;
        1078:  q   <=  32'b00000000000000000000000000000000 ;
        1079:  q   <=  32'b00000000000000000000000000000000 ;
        1080:  q   <=  32'b00000000000000000000000000000000 ;
        1081:  q   <=  32'b00000000000000000000000000000000 ;
        1082:  q   <=  32'b00000000000000000000000000000000 ;
        1083:  q   <=  32'b00000000000000000000000000000000 ;
        1084:  q   <=  32'b00000000000000000000000000000000 ;
        1085:  q   <=  32'b00000000000000000000000000000000 ;
        1086:  q   <=  32'b00000000000000000000000000000000 ;
        1087:  q   <=  32'b00000000000000000000000000000000 ;
        1088:  q   <=  32'b00000000000000000000000000000000 ;
        1089:  q   <=  32'b00000000000000000000000000000000 ;
        1090:  q   <=  32'b00000000000000000000000000000000 ;
        1091:  q   <=  32'b00000000000000000000000000000000 ;
        1092:  q   <=  32'b00000000000000000000000000000000 ;
        1093:  q   <=  32'b00000000000000000000000000000000 ;
        1094:  q   <=  32'b00000000000000000000000000000000 ;
        1095:  q   <=  32'b00000000000000000000000000000000 ;
        1096:  q   <=  32'b00000000000000000000000000000000 ;
        1097:  q   <=  32'b00000000000000000000000000000000 ;
        1098:  q   <=  32'b00000000000000000000000000000000 ;
        1099:  q   <=  32'b00000000000000000000000000000000 ;
        1100:  q   <=  32'b00000000000000000000000000000000 ;
        1101:  q   <=  32'b00000000000000000000000000000000 ;
        1102:  q   <=  32'b00000000000000000000000000000000 ;
        1103:  q   <=  32'b00000000000000000000000000000000 ;
        1104:  q   <=  32'b00000000000000000000000000000000 ;
        1105:  q   <=  32'b00000000000000000000000000000000 ;
        1106:  q   <=  32'b00000000000000000000000000000000 ;
        1107:  q   <=  32'b00000000000000000000000000000000 ;
        1108:  q   <=  32'b00000000000000000000000000000000 ;
        1109:  q   <=  32'b00000000000000000000000000000000 ;
        1110:  q   <=  32'b00000000000000000000000000000000 ;
        1111:  q   <=  32'b00000000000000000000000000000000 ;
        1112:  q   <=  32'b00000000000000000000000000000000 ;
        1113:  q   <=  32'b00000000000000000000000000000000 ;
        1114:  q   <=  32'b00000000000000000000000000000000 ;
        1115:  q   <=  32'b00000000000000000000000000000000 ;
        1116:  q   <=  32'b00000000000000000000000000000000 ;
        1117:  q   <=  32'b00000000000000000000000000000000 ;
        1118:  q   <=  32'b00000000000000000000000000000000 ;
        1119:  q   <=  32'b00000000000000000000000000000000 ;
        1120:  q   <=  32'b00000000000000000000000000000000 ;
        1121:  q   <=  32'b00000000000000000000000000000000 ;
        1122:  q   <=  32'b00000000000000000000000000000000 ;
        1123:  q   <=  32'b00000000000000000000000000000000 ;
        1124:  q   <=  32'b00000000000000000000000000000000 ;
        1125:  q   <=  32'b00000000000000000000000000000000 ;
        1126:  q   <=  32'b00000000000000000000000000000000 ;
        1127:  q   <=  32'b00000000000000000000000000000000 ;
        1128:  q   <=  32'b00000000000000000000000000000000 ;
        1129:  q   <=  32'b00000000000000000000000000000000 ;
        1130:  q   <=  32'b00000000000000000000000000000000 ;
        1131:  q   <=  32'b00000000000000000000000000000000 ;
        1132:  q   <=  32'b00000000000000000000000000000000 ;
        1133:  q   <=  32'b00000000000000000000000000000000 ;
        1134:  q   <=  32'b00000000000000000000000000000000 ;
        1135:  q   <=  32'b00000000000000000000000000000000 ;
        1136:  q   <=  32'b00000000000000000000000000000000 ;
        1137:  q   <=  32'b00000000000000000000000000000000 ;
        1138:  q   <=  32'b00000000000000000000000000000000 ;
        1139:  q   <=  32'b00000000000000000000000000000000 ;
        1140:  q   <=  32'b00000000000000000000000000000000 ;
        1141:  q   <=  32'b00000000000000000000000000000000 ;
        1142:  q   <=  32'b00000000000000000000000000000000 ;
        1143:  q   <=  32'b00000000000000000000000000000000 ;
        1144:  q   <=  32'b00000000000000000000000000000000 ;
        1145:  q   <=  32'b00000000000000000000000000000000 ;
        1146:  q   <=  32'b00000000000000000000000000000000 ;
        1147:  q   <=  32'b00000000000000000000000000000000 ;
        1148:  q   <=  32'b00000000000000000000000000000000 ;
        1149:  q   <=  32'b00000000000000000000000000000000 ;
        1150:  q   <=  32'b00000000000000000000000000000000 ;
        1151:  q   <=  32'b00000000000000000000000000000000 ;
        1152:  q   <=  32'b00000000000000000000000000000000 ;
        1153:  q   <=  32'b00000000000000000000000000000000 ;
        1154:  q   <=  32'b00000000000000000000000000000000 ;
        1155:  q   <=  32'b00000000000000000000000000000000 ;
        1156:  q   <=  32'b00000000000000000000000000000000 ;
        1157:  q   <=  32'b00000000000000000000000000000000 ;
        1158:  q   <=  32'b00000000000000000000000000000000 ;
        1159:  q   <=  32'b00000000000000000000000000000000 ;
        1160:  q   <=  32'b00000000000000000000000000000000 ;
        1161:  q   <=  32'b00000000000000000000000000000000 ;
        1162:  q   <=  32'b00000000000000000000000000000000 ;
        1163:  q   <=  32'b00000000000000000000000000000000 ;
        1164:  q   <=  32'b00000000000000000000000000000000 ;
        1165:  q   <=  32'b00000000000000000000000000000000 ;
        1166:  q   <=  32'b00000000000000000000000000000000 ;
        1167:  q   <=  32'b00000000000000000000000000000000 ;
        1168:  q   <=  32'b00000000000000000000000000000000 ;
        1169:  q   <=  32'b00000000000000000000000000000000 ;
        1170:  q   <=  32'b00000000000000000000000000000000 ;
        1171:  q   <=  32'b00000000000000000000000000000000 ;
        1172:  q   <=  32'b00000000000000000000000000000000 ;
        1173:  q   <=  32'b00000000000000000000000000000000 ;
        1174:  q   <=  32'b00000000000000000000000000000000 ;
        1175:  q   <=  32'b00000000000000000000000000000000 ;
        1176:  q   <=  32'b00000000000000000000000000000000 ;
        1177:  q   <=  32'b00111101110000011011100101011001 ;
        1178:  q   <=  32'b00111110110100101010001100001010 ;
        1179:  q   <=  32'b00111111001110011101011111001101 ;
        1180:  q   <=  32'b00111111100001001110010111001011 ;
        1181:  q   <=  32'b00111111101011001001011100111000 ;
        1182:  q   <=  32'b00111111110101000000000011110010 ;
        1183:  q   <=  32'b00111111111110110010001110111011 ;
        1184:  q   <=  32'b00111111110111011111111110101111 ;
        1185:  q   <=  32'b00111111101101110110100010010001 ;
        1186:  q   <=  32'b00111111100100010001011000101111 ;
        1187:  q   <=  32'b00111111010101100000111110101000 ;
        1188:  q   <=  32'b00111111000010100111100110010100 ;
        1189:  q   <=  32'b00111110011111011010001100000000 ;
        1190:  q   <=  32'b00000000000000000000000000000000 ;
        1191:  q   <=  32'b00000000000000000000000000000000 ;
        1192:  q   <=  32'b00000000000000000000000000000000 ;
        1193:  q   <=  32'b00000000000000000000000000000000 ;
        1194:  q   <=  32'b00000000000000000000000000000000 ;
        1195:  q   <=  32'b00000000000000000000000000000000 ;
        1196:  q   <=  32'b00000000000000000000000000000000 ;
        1197:  q   <=  32'b00000000000000000000000000000000 ;
        1198:  q   <=  32'b00000000000000000000000000000000 ;
        1199:  q   <=  32'b00000000000000000000000000000000 ;
        1200:  q   <=  32'b00000000000000000000000000000000 ;
        1201:  q   <=  32'b00000000000000000000000000000000 ;
        1202:  q   <=  32'b00000000000000000000000000000000 ;
        1203:  q   <=  32'b00000000000000000000000000000000 ;
        1204:  q   <=  32'b00000000000000000000000000000000 ;
        1205:  q   <=  32'b00000000000000000000000000000000 ;
        1206:  q   <=  32'b00000000000000000000000000000000 ;
        1207:  q   <=  32'b00000000000000000000000000000000 ;
        1208:  q   <=  32'b00000000000000000000000000000000 ;
        1209:  q   <=  32'b00000000000000000000000000000000 ;
        1210:  q   <=  32'b00000000000000000000000000000000 ;
        1211:  q   <=  32'b00000000000000000000000000000000 ;
        1212:  q   <=  32'b00000000000000000000000000000000 ;
        1213:  q   <=  32'b00000000000000000000000000000000 ;
        1214:  q   <=  32'b00000000000000000000000000000000 ;
        1215:  q   <=  32'b00000000000000000000000000000000 ;
        1216:  q   <=  32'b00000000000000000000000000000000 ;
        1217:  q   <=  32'b00000000000000000000000000000000 ;
        1218:  q   <=  32'b00000000000000000000000000000000 ;
        1219:  q   <=  32'b00000000000000000000000000000000 ;
        1220:  q   <=  32'b00000000000000000000000000000000 ;
        1221:  q   <=  32'b00000000000000000000000000000000 ;
        1222:  q   <=  32'b00000000000000000000000000000000 ;
        1223:  q   <=  32'b00000000000000000000000000000000 ;
        1224:  q   <=  32'b00000000000000000000000000000000 ;
        1225:  q   <=  32'b00000000000000000000000000000000 ;
        1226:  q   <=  32'b00000000000000000000000000000000 ;
        1227:  q   <=  32'b00000000000000000000000000000000 ;
        1228:  q   <=  32'b00000000000000000000000000000000 ;
        1229:  q   <=  32'b00000000000000000000000000000000 ;
        1230:  q   <=  32'b00000000000000000000000000000000 ;
        1231:  q   <=  32'b00000000000000000000000000000000 ;
        1232:  q   <=  32'b00000000000000000000000000000000 ;
        1233:  q   <=  32'b00000000000000000000000000000000 ;
        1234:  q   <=  32'b00000000000000000000000000000000 ;
        1235:  q   <=  32'b00000000000000000000000000000000 ;
        1236:  q   <=  32'b00000000000000000000000000000000 ;
        1237:  q   <=  32'b00000000000000000000000000000000 ;
        1238:  q   <=  32'b00000000000000000000000000000000 ;
        1239:  q   <=  32'b00000000000000000000000000000000 ;
        1240:  q   <=  32'b00000000000000000000000000000000 ;
        1241:  q   <=  32'b00000000000000000000000000000000 ;
        1242:  q   <=  32'b00000000000000000000000000000000 ;
        1243:  q   <=  32'b00000000000000000000000000000000 ;
        1244:  q   <=  32'b00000000000000000000000000000000 ;
        1245:  q   <=  32'b00000000000000000000000000000000 ;
        1246:  q   <=  32'b00000000000000000000000000000000 ;
        1247:  q   <=  32'b00000000000000000000000000000000 ;
        1248:  q   <=  32'b00000000000000000000000000000000 ;
        1249:  q   <=  32'b00000000000000000000000000000000 ;
        1250:  q   <=  32'b00000000000000000000000000000000 ;
        1251:  q   <=  32'b00000000000000000000000000000000 ;
        1252:  q   <=  32'b00000000000000000000000000000000 ;
        1253:  q   <=  32'b00000000000000000000000000000000 ;
        1254:  q   <=  32'b00000000000000000000000000000000 ;
        1255:  q   <=  32'b00000000000000000000000000000000 ;
        1256:  q   <=  32'b00000000000000000000000000000000 ;
        1257:  q   <=  32'b00000000000000000000000000000000 ;
        1258:  q   <=  32'b00000000000000000000000000000000 ;
        1259:  q   <=  32'b00000000000000000000000000000000 ;
        1260:  q   <=  32'b00000000000000000000000000000000 ;
        1261:  q   <=  32'b00000000000000000000000000000000 ;
        1262:  q   <=  32'b00000000000000000000000000000000 ;
        1263:  q   <=  32'b00000000000000000000000000000000 ;
        1264:  q   <=  32'b00000000000000000000000000000000 ;
        1265:  q   <=  32'b00000000000000000000000000000000 ;
        1266:  q   <=  32'b00000000000000000000000000000000 ;
        1267:  q   <=  32'b00000000000000000000000000000000 ;
        1268:  q   <=  32'b00000000000000000000000000000000 ;
        1269:  q   <=  32'b00000000000000000000000000000000 ;
        1270:  q   <=  32'b00000000000000000000000000000000 ;
        1271:  q   <=  32'b00000000000000000000000000000000 ;
        1272:  q   <=  32'b00000000000000000000000000000000 ;
        1273:  q   <=  32'b00000000000000000000000000000000 ;
        1274:  q   <=  32'b00000000000000000000000000000000 ;
        1275:  q   <=  32'b00000000000000000000000000000000 ;
        1276:  q   <=  32'b00000000000000000000000000000000 ;
        1277:  q   <=  32'b00000000000000000000000000000000 ;
        1278:  q   <=  32'b00000000000000000000000000000000 ;
        1279:  q   <=  32'b00000000000000000000000000000000 ;
        1280:  q   <=  32'b00000000000000000000000000000000 ;
        1281:  q   <=  32'b00000000000000000000000000000000 ;
        1282:  q   <=  32'b00000000000000000000000000000000 ;
        1283:  q   <=  32'b00000000000000000000000000000000 ;
        1284:  q   <=  32'b00000000000000000000000000000000 ;
        1285:  q   <=  32'b00000000000000000000000000000000 ;
        1286:  q   <=  32'b00000000000000000000000000000000 ;
        1287:  q   <=  32'b00000000000000000000000000000000 ;
        1288:  q   <=  32'b00000000000000000000000000000000 ;
        1289:  q   <=  32'b00000000000000000000000000000000 ;
        1290:  q   <=  32'b00000000000000000000000000000000 ;
        1291:  q   <=  32'b00000000000000000000000000000000 ;
        1292:  q   <=  32'b00000000000000000000000000000000 ;
        1293:  q   <=  32'b00000000000000000000000000000000 ;
        1294:  q   <=  32'b00000000000000000000000000000000 ;
        1295:  q   <=  32'b00000000000000000000000000000000 ;
        1296:  q   <=  32'b00000000000000000000000000000000 ;
        1297:  q   <=  32'b00000000000000000000000000000000 ;
        1298:  q   <=  32'b00000000000000000000000000000000 ;
        1299:  q   <=  32'b00000000000000000000000000000000 ;
        1300:  q   <=  32'b00000000000000000000000000000000 ;
        1301:  q   <=  32'b00000000000000000000000000000000 ;
        1302:  q   <=  32'b00000000000000000000000000000000 ;
        1303:  q   <=  32'b00000000000000000000000000000000 ;
        1304:  q   <=  32'b00000000000000000000000000000000 ;
        1305:  q   <=  32'b00000000000000000000000000000000 ;
        1306:  q   <=  32'b00000000000000000000000000000000 ;
        1307:  q   <=  32'b00000000000000000000000000000000 ;
        1308:  q   <=  32'b00000000000000000000000000000000 ;
        1309:  q   <=  32'b00000000000000000000000000000000 ;
        1310:  q   <=  32'b00000000000000000000000000000000 ;
        1311:  q   <=  32'b00000000000000000000000000000000 ;
        1312:  q   <=  32'b00000000000000000000000000000000 ;
        1313:  q   <=  32'b00000000000000000000000000000000 ;
        1314:  q   <=  32'b00000000000000000000000000000000 ;
        1315:  q   <=  32'b00000000000000000000000000000000 ;
        1316:  q   <=  32'b00000000000000000000000000000000 ;
        1317:  q   <=  32'b00000000000000000000000000000000 ;
        1318:  q   <=  32'b00000000000000000000000000000000 ;
        1319:  q   <=  32'b00000000000000000000000000000000 ;
        1320:  q   <=  32'b00000000000000000000000000000000 ;
        1321:  q   <=  32'b00000000000000000000000000000000 ;
        1322:  q   <=  32'b00000000000000000000000000000000 ;
        1323:  q   <=  32'b00000000000000000000000000000000 ;
        1324:  q   <=  32'b00000000000000000000000000000000 ;
        1325:  q   <=  32'b00000000000000000000000000000000 ;
        1326:  q   <=  32'b00000000000000000000000000000000 ;
        1327:  q   <=  32'b00000000000000000000000000000000 ;
        1328:  q   <=  32'b00000000000000000000000000000000 ;
        1329:  q   <=  32'b00000000000000000000000000000000 ;
        1330:  q   <=  32'b00000000000000000000000000000000 ;
        1331:  q   <=  32'b00000000000000000000000000000000 ;
        1332:  q   <=  32'b00000000000000000000000000000000 ;
        1333:  q   <=  32'b00000000000000000000000000000000 ;
        1334:  q   <=  32'b00000000000000000000000000000000 ;
        1335:  q   <=  32'b00000000000000000000000000000000 ;
        1336:  q   <=  32'b00000000000000000000000000000000 ;
        1337:  q   <=  32'b00000000000000000000000000000000 ;
        1338:  q   <=  32'b00000000000000000000000000000000 ;
        1339:  q   <=  32'b00000000000000000000000000000000 ;
        1340:  q   <=  32'b00000000000000000000000000000000 ;
        1341:  q   <=  32'b00000000000000000000000000000000 ;
        1342:  q   <=  32'b00000000000000000000000000000000 ;
        1343:  q   <=  32'b00000000000000000000000000000000 ;
        1344:  q   <=  32'b00000000000000000000000000000000 ;
        1345:  q   <=  32'b00000000000000000000000000000000 ;
        1346:  q   <=  32'b00000000000000000000000000000000 ;
        1347:  q   <=  32'b00000000000000000000000000000000 ;
        1348:  q   <=  32'b00000000000000000000000000000000 ;
        1349:  q   <=  32'b00000000000000000000000000000000 ;
        1350:  q   <=  32'b00000000000000000000000000000000 ;
        1351:  q   <=  32'b00000000000000000000000000000000 ;
        1352:  q   <=  32'b00000000000000000000000000000000 ;
        1353:  q   <=  32'b00000000000000000000000000000000 ;
        1354:  q   <=  32'b00000000000000000000000000000000 ;
        1355:  q   <=  32'b00000000000000000000000000000000 ;
        1356:  q   <=  32'b00000000000000000000000000000000 ;
        1357:  q   <=  32'b00000000000000000000000000000000 ;
        1358:  q   <=  32'b00000000000000000000000000000000 ;
        1359:  q   <=  32'b00000000000000000000000000000000 ;
        1360:  q   <=  32'b00000000000000000000000000000000 ;
        1361:  q   <=  32'b00000000000000000000000000000000 ;
        1362:  q   <=  32'b00000000000000000000000000000000 ;
        1363:  q   <=  32'b00000000000000000000000000000000 ;
        1364:  q   <=  32'b00000000000000000000000000000000 ;
        1365:  q   <=  32'b00000000000000000000000000000000 ;
        1366:  q   <=  32'b00000000000000000000000000000000 ;
        1367:  q   <=  32'b00000000000000000000000000000000 ;
        1368:  q   <=  32'b00000000000000000000000000000000 ;
        1369:  q   <=  32'b00000000000000000000000000000000 ;
        1370:  q   <=  32'b00000000000000000000000000000000 ;
        1371:  q   <=  32'b00000000000000000000000000000000 ;
        1372:  q   <=  32'b00000000000000000000000000000000 ;
        1373:  q   <=  32'b00000000000000000000000000000000 ;
        1374:  q   <=  32'b00000000000000000000000000000000 ;
        1375:  q   <=  32'b00000000000000000000000000000000 ;
        1376:  q   <=  32'b00000000000000000000000000000000 ;
        1377:  q   <=  32'b00000000000000000000000000000000 ;
        1378:  q   <=  32'b00000000000000000000000000000000 ;
        1379:  q   <=  32'b00000000000000000000000000000000 ;
        1380:  q   <=  32'b00000000000000000000000000000000 ;
        1381:  q   <=  32'b00000000000000000000000000000000 ;
        1382:  q   <=  32'b00000000000000000000000000000000 ;
        1383:  q   <=  32'b00000000000000000000000000000000 ;
        1384:  q   <=  32'b00000000000000000000000000000000 ;
        1385:  q   <=  32'b00000000000000000000000000000000 ;
        1386:  q   <=  32'b00000000000000000000000000000000 ;
        1387:  q   <=  32'b00000000000000000000000000000000 ;
        1388:  q   <=  32'b00000000000000000000000000000000 ;
        1389:  q   <=  32'b00000000000000000000000000000000 ;
        1390:  q   <=  32'b00000000000000000000000000000000 ;
        1391:  q   <=  32'b00000000000000000000000000000000 ;
        1392:  q   <=  32'b00000000000000000000000000000000 ;
        1393:  q   <=  32'b00000000000000000000000000000000 ;
        1394:  q   <=  32'b00000000000000000000000000000000 ;
        1395:  q   <=  32'b00000000000000000000000000000000 ;
        1396:  q   <=  32'b00000000000000000000000000000000 ;
        1397:  q   <=  32'b00000000000000000000000000000000 ;
        1398:  q   <=  32'b00000000000000000000000000000000 ;
        1399:  q   <=  32'b00000000000000000000000000000000 ;
        1400:  q   <=  32'b00000000000000000000000000000000 ;
        1401:  q   <=  32'b00000000000000000000000000000000 ;
        1402:  q   <=  32'b00000000000000000000000000000000 ;
        1403:  q   <=  32'b00000000000000000000000000000000 ;
        1404:  q   <=  32'b00000000000000000000000000000000 ;
        1405:  q   <=  32'b00000000000000000000000000000000 ;
        1406:  q   <=  32'b00000000000000000000000000000000 ;
        1407:  q   <=  32'b00000000000000000000000000000000 ;
        1408:  q   <=  32'b00000000000000000000000000000000 ;
        1409:  q   <=  32'b00000000000000000000000000000000 ;
        1410:  q   <=  32'b00000000000000000000000000000000 ;
        1411:  q   <=  32'b00000000000000000000000000000000 ;
        1412:  q   <=  32'b00000000000000000000000000000000 ;
        1413:  q   <=  32'b00000000000000000000000000000000 ;
        1414:  q   <=  32'b00000000000000000000000000000000 ;
        1415:  q   <=  32'b00000000000000000000000000000000 ;
        1416:  q   <=  32'b00000000000000000000000000000000 ;
        1417:  q   <=  32'b00000000000000000000000000000000 ;
        1418:  q   <=  32'b00000000000000000000000000000000 ;
        1419:  q   <=  32'b00000000000000000000000000000000 ;
        1420:  q   <=  32'b00000000000000000000000000000000 ;
        1421:  q   <=  32'b00000000000000000000000000000000 ;
        1422:  q   <=  32'b00000000000000000000000000000000 ;
        1423:  q   <=  32'b00000000000000000000000000000000 ;
        1424:  q   <=  32'b00000000000000000000000000000000 ;
        1425:  q   <=  32'b00000000000000000000000000000000 ;
        1426:  q   <=  32'b00000000000000000000000000000000 ;
        1427:  q   <=  32'b00000000000000000000000000000000 ;
        1428:  q   <=  32'b00000000000000000000000000000000 ;
        1429:  q   <=  32'b00000000000000000000000000000000 ;
        1430:  q   <=  32'b00000000000000000000000000000000 ;
        1431:  q   <=  32'b00000000000000000000000000000000 ;
        1432:  q   <=  32'b00000000000000000000000000000000 ;
        1433:  q   <=  32'b00000000000000000000000000000000 ;
        1434:  q   <=  32'b00000000000000000000000000000000 ;
        1435:  q   <=  32'b00000000000000000000000000000000 ;
        1436:  q   <=  32'b00000000000000000000000000000000 ;
        1437:  q   <=  32'b00000000000000000000000000000000 ;
        1438:  q   <=  32'b00000000000000000000000000000000 ;
        1439:  q   <=  32'b00000000000000000000000000000000 ;
        1440:  q   <=  32'b00111110100010000000000101000001 ;
        1441:  q   <=  32'b00111111000100010010111011011101 ;
        1442:  q   <=  32'b00111111010111011101001110100000 ;
        1443:  q   <=  32'b00111111100101001111100000101011 ;
        1444:  q   <=  32'b00111111101110101100001100110101 ;
        1445:  q   <=  32'b00111111111000000100101110011111 ;
        1446:  q   <=  32'b00111111111110100110110111100101 ;
        1447:  q   <=  32'b00111111110101010110100010101110 ;
        1448:  q   <=  32'b00111111101100001010010000001111 ;
        1449:  q   <=  32'b00111111100011000001111101011111 ;
        1450:  q   <=  32'b00111111010011111011001111110001 ;
        1451:  q   <=  32'b00111111000001111010011001101111 ;
        1452:  q   <=  32'b00111110100000000010100111101001 ;
        1453:  q   <=  32'b00000000000000000000000000000000 ;
        1454:  q   <=  32'b00000000000000000000000000000000 ;
        1455:  q   <=  32'b00000000000000000000000000000000 ;
        1456:  q   <=  32'b00000000000000000000000000000000 ;
        1457:  q   <=  32'b00000000000000000000000000000000 ;
        1458:  q   <=  32'b00000000000000000000000000000000 ;
        1459:  q   <=  32'b00000000000000000000000000000000 ;
        1460:  q   <=  32'b00000000000000000000000000000000 ;
        1461:  q   <=  32'b00000000000000000000000000000000 ;
        1462:  q   <=  32'b00000000000000000000000000000000 ;
        1463:  q   <=  32'b00000000000000000000000000000000 ;
        1464:  q   <=  32'b00000000000000000000000000000000 ;
        1465:  q   <=  32'b00000000000000000000000000000000 ;
        1466:  q   <=  32'b00000000000000000000000000000000 ;
        1467:  q   <=  32'b00000000000000000000000000000000 ;
        1468:  q   <=  32'b00000000000000000000000000000000 ;
        1469:  q   <=  32'b00000000000000000000000000000000 ;
        1470:  q   <=  32'b00000000000000000000000000000000 ;
        1471:  q   <=  32'b00000000000000000000000000000000 ;
        1472:  q   <=  32'b00000000000000000000000000000000 ;
        1473:  q   <=  32'b00000000000000000000000000000000 ;
        1474:  q   <=  32'b00000000000000000000000000000000 ;
        1475:  q   <=  32'b00000000000000000000000000000000 ;
        1476:  q   <=  32'b00000000000000000000000000000000 ;
        1477:  q   <=  32'b00000000000000000000000000000000 ;
        1478:  q   <=  32'b00000000000000000000000000000000 ;
        1479:  q   <=  32'b00000000000000000000000000000000 ;
        1480:  q   <=  32'b00000000000000000000000000000000 ;
        1481:  q   <=  32'b00000000000000000000000000000000 ;
        1482:  q   <=  32'b00000000000000000000000000000000 ;
        1483:  q   <=  32'b00000000000000000000000000000000 ;
        1484:  q   <=  32'b00000000000000000000000000000000 ;
        1485:  q   <=  32'b00000000000000000000000000000000 ;
        1486:  q   <=  32'b00000000000000000000000000000000 ;
        1487:  q   <=  32'b00000000000000000000000000000000 ;
        1488:  q   <=  32'b00000000000000000000000000000000 ;
        1489:  q   <=  32'b00000000000000000000000000000000 ;
        1490:  q   <=  32'b00000000000000000000000000000000 ;
        1491:  q   <=  32'b00000000000000000000000000000000 ;
        1492:  q   <=  32'b00000000000000000000000000000000 ;
        1493:  q   <=  32'b00000000000000000000000000000000 ;
        1494:  q   <=  32'b00000000000000000000000000000000 ;
        1495:  q   <=  32'b00000000000000000000000000000000 ;
        1496:  q   <=  32'b00000000000000000000000000000000 ;
        1497:  q   <=  32'b00000000000000000000000000000000 ;
        1498:  q   <=  32'b00000000000000000000000000000000 ;
        1499:  q   <=  32'b00000000000000000000000000000000 ;
        1500:  q   <=  32'b00000000000000000000000000000000 ;
        1501:  q   <=  32'b00000000000000000000000000000000 ;
        1502:  q   <=  32'b00000000000000000000000000000000 ;
        1503:  q   <=  32'b00000000000000000000000000000000 ;
        1504:  q   <=  32'b00000000000000000000000000000000 ;
        1505:  q   <=  32'b00000000000000000000000000000000 ;
        1506:  q   <=  32'b00000000000000000000000000000000 ;
        1507:  q   <=  32'b00000000000000000000000000000000 ;
        1508:  q   <=  32'b00000000000000000000000000000000 ;
        1509:  q   <=  32'b00000000000000000000000000000000 ;
        1510:  q   <=  32'b00000000000000000000000000000000 ;
        1511:  q   <=  32'b00000000000000000000000000000000 ;
        1512:  q   <=  32'b00000000000000000000000000000000 ;
        1513:  q   <=  32'b00000000000000000000000000000000 ;
        1514:  q   <=  32'b00000000000000000000000000000000 ;
        1515:  q   <=  32'b00000000000000000000000000000000 ;
        1516:  q   <=  32'b00000000000000000000000000000000 ;
        1517:  q   <=  32'b00000000000000000000000000000000 ;
        1518:  q   <=  32'b00000000000000000000000000000000 ;
        1519:  q   <=  32'b00000000000000000000000000000000 ;
        1520:  q   <=  32'b00000000000000000000000000000000 ;
        1521:  q   <=  32'b00000000000000000000000000000000 ;
        1522:  q   <=  32'b00000000000000000000000000000000 ;
        1523:  q   <=  32'b00000000000000000000000000000000 ;
        1524:  q   <=  32'b00000000000000000000000000000000 ;
        1525:  q   <=  32'b00000000000000000000000000000000 ;
        1526:  q   <=  32'b00000000000000000000000000000000 ;
        1527:  q   <=  32'b00000000000000000000000000000000 ;
        1528:  q   <=  32'b00000000000000000000000000000000 ;
        1529:  q   <=  32'b00000000000000000000000000000000 ;
        1530:  q   <=  32'b00000000000000000000000000000000 ;
        1531:  q   <=  32'b00000000000000000000000000000000 ;
        1532:  q   <=  32'b00000000000000000000000000000000 ;
        1533:  q   <=  32'b00000000000000000000000000000000 ;
        1534:  q   <=  32'b00000000000000000000000000000000 ;
        1535:  q   <=  32'b00000000000000000000000000000000 ;
        1536:  q   <=  32'b00000000000000000000000000000000 ;
        1537:  q   <=  32'b00000000000000000000000000000000 ;
        1538:  q   <=  32'b00000000000000000000000000000000 ;
        1539:  q   <=  32'b00000000000000000000000000000000 ;
        1540:  q   <=  32'b00000000000000000000000000000000 ;
        1541:  q   <=  32'b00000000000000000000000000000000 ;
        1542:  q   <=  32'b00000000000000000000000000000000 ;
        1543:  q   <=  32'b00000000000000000000000000000000 ;
        1544:  q   <=  32'b00000000000000000000000000000000 ;
        1545:  q   <=  32'b00000000000000000000000000000000 ;
        1546:  q   <=  32'b00000000000000000000000000000000 ;
        1547:  q   <=  32'b00000000000000000000000000000000 ;
        1548:  q   <=  32'b00000000000000000000000000000000 ;
        1549:  q   <=  32'b00000000000000000000000000000000 ;
        1550:  q   <=  32'b00000000000000000000000000000000 ;
        1551:  q   <=  32'b00000000000000000000000000000000 ;
        1552:  q   <=  32'b00000000000000000000000000000000 ;
        1553:  q   <=  32'b00000000000000000000000000000000 ;
        1554:  q   <=  32'b00000000000000000000000000000000 ;
        1555:  q   <=  32'b00000000000000000000000000000000 ;
        1556:  q   <=  32'b00000000000000000000000000000000 ;
        1557:  q   <=  32'b00000000000000000000000000000000 ;
        1558:  q   <=  32'b00000000000000000000000000000000 ;
        1559:  q   <=  32'b00000000000000000000000000000000 ;
        1560:  q   <=  32'b00000000000000000000000000000000 ;
        1561:  q   <=  32'b00000000000000000000000000000000 ;
        1562:  q   <=  32'b00000000000000000000000000000000 ;
        1563:  q   <=  32'b00000000000000000000000000000000 ;
        1564:  q   <=  32'b00000000000000000000000000000000 ;
        1565:  q   <=  32'b00000000000000000000000000000000 ;
        1566:  q   <=  32'b00000000000000000000000000000000 ;
        1567:  q   <=  32'b00000000000000000000000000000000 ;
        1568:  q   <=  32'b00000000000000000000000000000000 ;
        1569:  q   <=  32'b00000000000000000000000000000000 ;
        1570:  q   <=  32'b00000000000000000000000000000000 ;
        1571:  q   <=  32'b00000000000000000000000000000000 ;
        1572:  q   <=  32'b00000000000000000000000000000000 ;
        1573:  q   <=  32'b00000000000000000000000000000000 ;
        1574:  q   <=  32'b00000000000000000000000000000000 ;
        1575:  q   <=  32'b00000000000000000000000000000000 ;
        1576:  q   <=  32'b00000000000000000000000000000000 ;
        1577:  q   <=  32'b00000000000000000000000000000000 ;
        1578:  q   <=  32'b00000000000000000000000000000000 ;
        1579:  q   <=  32'b00000000000000000000000000000000 ;
        1580:  q   <=  32'b00000000000000000000000000000000 ;
        1581:  q   <=  32'b00000000000000000000000000000000 ;
        1582:  q   <=  32'b00000000000000000000000000000000 ;
        1583:  q   <=  32'b00000000000000000000000000000000 ;
        1584:  q   <=  32'b00000000000000000000000000000000 ;
        1585:  q   <=  32'b00000000000000000000000000000000 ;
        1586:  q   <=  32'b00000000000000000000000000000000 ;
        1587:  q   <=  32'b00000000000000000000000000000000 ;
        1588:  q   <=  32'b00000000000000000000000000000000 ;
        1589:  q   <=  32'b00000000000000000000000000000000 ;
        1590:  q   <=  32'b00000000000000000000000000000000 ;
        1591:  q   <=  32'b00000000000000000000000000000000 ;
        1592:  q   <=  32'b00000000000000000000000000000000 ;
        1593:  q   <=  32'b00000000000000000000000000000000 ;
        1594:  q   <=  32'b00000000000000000000000000000000 ;
        1595:  q   <=  32'b00000000000000000000000000000000 ;
        1596:  q   <=  32'b00000000000000000000000000000000 ;
        1597:  q   <=  32'b00000000000000000000000000000000 ;
        1598:  q   <=  32'b00000000000000000000000000000000 ;
        1599:  q   <=  32'b00000000000000000000000000000000 ;
        1600:  q   <=  32'b00000000000000000000000000000000 ;
        1601:  q   <=  32'b00000000000000000000000000000000 ;
        1602:  q   <=  32'b00000000000000000000000000000000 ;
        1603:  q   <=  32'b00000000000000000000000000000000 ;
        1604:  q   <=  32'b00000000000000000000000000000000 ;
        1605:  q   <=  32'b00000000000000000000000000000000 ;
        1606:  q   <=  32'b00000000000000000000000000000000 ;
        1607:  q   <=  32'b00000000000000000000000000000000 ;
        1608:  q   <=  32'b00000000000000000000000000000000 ;
        1609:  q   <=  32'b00000000000000000000000000000000 ;
        1610:  q   <=  32'b00000000000000000000000000000000 ;
        1611:  q   <=  32'b00000000000000000000000000000000 ;
        1612:  q   <=  32'b00000000000000000000000000000000 ;
        1613:  q   <=  32'b00000000000000000000000000000000 ;
        1614:  q   <=  32'b00000000000000000000000000000000 ;
        1615:  q   <=  32'b00000000000000000000000000000000 ;
        1616:  q   <=  32'b00000000000000000000000000000000 ;
        1617:  q   <=  32'b00000000000000000000000000000000 ;
        1618:  q   <=  32'b00000000000000000000000000000000 ;
        1619:  q   <=  32'b00000000000000000000000000000000 ;
        1620:  q   <=  32'b00000000000000000000000000000000 ;
        1621:  q   <=  32'b00000000000000000000000000000000 ;
        1622:  q   <=  32'b00000000000000000000000000000000 ;
        1623:  q   <=  32'b00000000000000000000000000000000 ;
        1624:  q   <=  32'b00000000000000000000000000000000 ;
        1625:  q   <=  32'b00000000000000000000000000000000 ;
        1626:  q   <=  32'b00000000000000000000000000000000 ;
        1627:  q   <=  32'b00000000000000000000000000000000 ;
        1628:  q   <=  32'b00000000000000000000000000000000 ;
        1629:  q   <=  32'b00000000000000000000000000000000 ;
        1630:  q   <=  32'b00000000000000000000000000000000 ;
        1631:  q   <=  32'b00000000000000000000000000000000 ;
        1632:  q   <=  32'b00000000000000000000000000000000 ;
        1633:  q   <=  32'b00000000000000000000000000000000 ;
        1634:  q   <=  32'b00000000000000000000000000000000 ;
        1635:  q   <=  32'b00000000000000000000000000000000 ;
        1636:  q   <=  32'b00000000000000000000000000000000 ;
        1637:  q   <=  32'b00000000000000000000000000000000 ;
        1638:  q   <=  32'b00000000000000000000000000000000 ;
        1639:  q   <=  32'b00000000000000000000000000000000 ;
        1640:  q   <=  32'b00000000000000000000000000000000 ;
        1641:  q   <=  32'b00000000000000000000000000000000 ;
        1642:  q   <=  32'b00000000000000000000000000000000 ;
        1643:  q   <=  32'b00000000000000000000000000000000 ;
        1644:  q   <=  32'b00000000000000000000000000000000 ;
        1645:  q   <=  32'b00000000000000000000000000000000 ;
        1646:  q   <=  32'b00000000000000000000000000000000 ;
        1647:  q   <=  32'b00000000000000000000000000000000 ;
        1648:  q   <=  32'b00000000000000000000000000000000 ;
        1649:  q   <=  32'b00000000000000000000000000000000 ;
        1650:  q   <=  32'b00000000000000000000000000000000 ;
        1651:  q   <=  32'b00000000000000000000000000000000 ;
        1652:  q   <=  32'b00000000000000000000000000000000 ;
        1653:  q   <=  32'b00000000000000000000000000000000 ;
        1654:  q   <=  32'b00000000000000000000000000000000 ;
        1655:  q   <=  32'b00000000000000000000000000000000 ;
        1656:  q   <=  32'b00000000000000000000000000000000 ;
        1657:  q   <=  32'b00000000000000000000000000000000 ;
        1658:  q   <=  32'b00000000000000000000000000000000 ;
        1659:  q   <=  32'b00000000000000000000000000000000 ;
        1660:  q   <=  32'b00000000000000000000000000000000 ;
        1661:  q   <=  32'b00000000000000000000000000000000 ;
        1662:  q   <=  32'b00000000000000000000000000000000 ;
        1663:  q   <=  32'b00000000000000000000000000000000 ;
        1664:  q   <=  32'b00000000000000000000000000000000 ;
        1665:  q   <=  32'b00000000000000000000000000000000 ;
        1666:  q   <=  32'b00000000000000000000000000000000 ;
        1667:  q   <=  32'b00000000000000000000000000000000 ;
        1668:  q   <=  32'b00000000000000000000000000000000 ;
        1669:  q   <=  32'b00000000000000000000000000000000 ;
        1670:  q   <=  32'b00000000000000000000000000000000 ;
        1671:  q   <=  32'b00000000000000000000000000000000 ;
        1672:  q   <=  32'b00000000000000000000000000000000 ;
        1673:  q   <=  32'b00000000000000000000000000000000 ;
        1674:  q   <=  32'b00000000000000000000000000000000 ;
        1675:  q   <=  32'b00000000000000000000000000000000 ;
        1676:  q   <=  32'b00000000000000000000000000000000 ;
        1677:  q   <=  32'b00000000000000000000000000000000 ;
        1678:  q   <=  32'b00000000000000000000000000000000 ;
        1679:  q   <=  32'b00000000000000000000000000000000 ;
        1680:  q   <=  32'b00000000000000000000000000000000 ;
        1681:  q   <=  32'b00000000000000000000000000000000 ;
        1682:  q   <=  32'b00000000000000000000000000000000 ;
        1683:  q   <=  32'b00000000000000000000000000000000 ;
        1684:  q   <=  32'b00000000000000000000000000000000 ;
        1685:  q   <=  32'b00000000000000000000000000000000 ;
        1686:  q   <=  32'b00000000000000000000000000000000 ;
        1687:  q   <=  32'b00000000000000000000000000000000 ;
        1688:  q   <=  32'b00000000000000000000000000000000 ;
        1689:  q   <=  32'b00000000000000000000000000000000 ;
        1690:  q   <=  32'b00000000000000000000000000000000 ;
        1691:  q   <=  32'b00000000000000000000000000000000 ;
        1692:  q   <=  32'b00000000000000000000000000000000 ;
        1693:  q   <=  32'b00000000000000000000000000000000 ;
        1694:  q   <=  32'b00000000000000000000000000000000 ;
        1695:  q   <=  32'b00000000000000000000000000000000 ;
        1696:  q   <=  32'b00000000000000000000000000000000 ;
        1697:  q   <=  32'b00000000000000000000000000000000 ;
        1698:  q   <=  32'b00000000000000000000000000000000 ;
        1699:  q   <=  32'b00000000000000000000000000000000 ;
        1700:  q   <=  32'b00000000000000000000000000000000 ;
        1701:  q   <=  32'b00000000000000000000000000000000 ;
        1702:  q   <=  32'b00111101001100100100001101000100 ;
        1703:  q   <=  32'b00111110101010100101110101000110 ;
        1704:  q   <=  32'b00111111000111101011011111100001 ;
        1705:  q   <=  32'b00111111011001111100000101000001 ;
        1706:  q   <=  32'b00111111100110000010011000000111 ;
        1707:  q   <=  32'b00111111101111000010110011001000 ;
        1708:  q   <=  32'b00111111110111111111010110000101 ;
        1709:  q   <=  32'b00111111111111000111111100100000 ;
        1710:  q   <=  32'b00111111110110010011000010001110 ;
        1711:  q   <=  32'b00111111101101100001111000100110 ;
        1712:  q   <=  32'b00111111100100110100011101010000 ;
        1713:  q   <=  32'b00111111011000010101011011101100 ;
        1714:  q   <=  32'b00111111000111001001010000000001 ;
        1715:  q   <=  32'b00111110101100001000100101110100 ;
        1716:  q   <=  32'b00111101101000110011111110100101 ;
        1717:  q   <=  32'b00000000000000000000000000000000 ;
        1718:  q   <=  32'b00000000000000000000000000000000 ;
        1719:  q   <=  32'b00000000000000000000000000000000 ;
        1720:  q   <=  32'b00000000000000000000000000000000 ;
        1721:  q   <=  32'b00000000000000000000000000000000 ;
        1722:  q   <=  32'b00000000000000000000000000000000 ;
        1723:  q   <=  32'b00000000000000000000000000000000 ;
        1724:  q   <=  32'b00000000000000000000000000000000 ;
        1725:  q   <=  32'b00000000000000000000000000000000 ;
        1726:  q   <=  32'b00000000000000000000000000000000 ;
        1727:  q   <=  32'b00000000000000000000000000000000 ;
        1728:  q   <=  32'b00000000000000000000000000000000 ;
        1729:  q   <=  32'b00000000000000000000000000000000 ;
        1730:  q   <=  32'b00000000000000000000000000000000 ;
        1731:  q   <=  32'b00000000000000000000000000000000 ;
        1732:  q   <=  32'b00000000000000000000000000000000 ;
        1733:  q   <=  32'b00000000000000000000000000000000 ;
        1734:  q   <=  32'b00000000000000000000000000000000 ;
        1735:  q   <=  32'b00000000000000000000000000000000 ;
        1736:  q   <=  32'b00000000000000000000000000000000 ;
        1737:  q   <=  32'b00000000000000000000000000000000 ;
        1738:  q   <=  32'b00000000000000000000000000000000 ;
        1739:  q   <=  32'b00000000000000000000000000000000 ;
        1740:  q   <=  32'b00000000000000000000000000000000 ;
        1741:  q   <=  32'b00000000000000000000000000000000 ;
        1742:  q   <=  32'b00000000000000000000000000000000 ;
        1743:  q   <=  32'b00000000000000000000000000000000 ;
        1744:  q   <=  32'b00000000000000000000000000000000 ;
        1745:  q   <=  32'b00000000000000000000000000000000 ;
        1746:  q   <=  32'b00000000000000000000000000000000 ;
        1747:  q   <=  32'b00000000000000000000000000000000 ;
        1748:  q   <=  32'b00000000000000000000000000000000 ;
        1749:  q   <=  32'b00000000000000000000000000000000 ;
        1750:  q   <=  32'b00000000000000000000000000000000 ;
        1751:  q   <=  32'b00000000000000000000000000000000 ;
        1752:  q   <=  32'b00000000000000000000000000000000 ;
        1753:  q   <=  32'b00000000000000000000000000000000 ;
        1754:  q   <=  32'b00000000000000000000000000000000 ;
        1755:  q   <=  32'b00000000000000000000000000000000 ;
        1756:  q   <=  32'b00000000000000000000000000000000 ;
        1757:  q   <=  32'b00000000000000000000000000000000 ;
        1758:  q   <=  32'b00000000000000000000000000000000 ;
        1759:  q   <=  32'b00000000000000000000000000000000 ;
        1760:  q   <=  32'b00000000000000000000000000000000 ;
        1761:  q   <=  32'b00000000000000000000000000000000 ;
        1762:  q   <=  32'b00000000000000000000000000000000 ;
        1763:  q   <=  32'b00000000000000000000000000000000 ;
        1764:  q   <=  32'b00000000000000000000000000000000 ;
        1765:  q   <=  32'b00000000000000000000000000000000 ;
        1766:  q   <=  32'b00000000000000000000000000000000 ;
        1767:  q   <=  32'b00000000000000000000000000000000 ;
        1768:  q   <=  32'b00000000000000000000000000000000 ;
        1769:  q   <=  32'b00000000000000000000000000000000 ;
        1770:  q   <=  32'b00000000000000000000000000000000 ;
        1771:  q   <=  32'b00000000000000000000000000000000 ;
        1772:  q   <=  32'b00000000000000000000000000000000 ;
        1773:  q   <=  32'b00000000000000000000000000000000 ;
        1774:  q   <=  32'b00000000000000000000000000000000 ;
        1775:  q   <=  32'b00000000000000000000000000000000 ;
        1776:  q   <=  32'b00000000000000000000000000000000 ;
        1777:  q   <=  32'b00000000000000000000000000000000 ;
        1778:  q   <=  32'b00000000000000000000000000000000 ;
        1779:  q   <=  32'b00000000000000000000000000000000 ;
        1780:  q   <=  32'b00000000000000000000000000000000 ;
        1781:  q   <=  32'b00000000000000000000000000000000 ;
        1782:  q   <=  32'b00000000000000000000000000000000 ;
        1783:  q   <=  32'b00000000000000000000000000000000 ;
        1784:  q   <=  32'b00000000000000000000000000000000 ;
        1785:  q   <=  32'b00000000000000000000000000000000 ;
        1786:  q   <=  32'b00000000000000000000000000000000 ;
        1787:  q   <=  32'b00000000000000000000000000000000 ;
        1788:  q   <=  32'b00000000000000000000000000000000 ;
        1789:  q   <=  32'b00000000000000000000000000000000 ;
        1790:  q   <=  32'b00000000000000000000000000000000 ;
        1791:  q   <=  32'b00000000000000000000000000000000 ;
        1792:  q   <=  32'b00000000000000000000000000000000 ;
        1793:  q   <=  32'b00000000000000000000000000000000 ;
        1794:  q   <=  32'b00000000000000000000000000000000 ;
        1795:  q   <=  32'b00000000000000000000000000000000 ;
        1796:  q   <=  32'b00000000000000000000000000000000 ;
        1797:  q   <=  32'b00000000000000000000000000000000 ;
        1798:  q   <=  32'b00000000000000000000000000000000 ;
        1799:  q   <=  32'b00000000000000000000000000000000 ;
        1800:  q   <=  32'b00000000000000000000000000000000 ;
        1801:  q   <=  32'b00000000000000000000000000000000 ;
        1802:  q   <=  32'b00000000000000000000000000000000 ;
        1803:  q   <=  32'b00000000000000000000000000000000 ;
        1804:  q   <=  32'b00000000000000000000000000000000 ;
        1805:  q   <=  32'b00000000000000000000000000000000 ;
        1806:  q   <=  32'b00000000000000000000000000000000 ;
        1807:  q   <=  32'b00000000000000000000000000000000 ;
        1808:  q   <=  32'b00000000000000000000000000000000 ;
        1809:  q   <=  32'b00000000000000000000000000000000 ;
        1810:  q   <=  32'b00000000000000000000000000000000 ;
        1811:  q   <=  32'b00000000000000000000000000000000 ;
        1812:  q   <=  32'b00000000000000000000000000000000 ;
        1813:  q   <=  32'b00000000000000000000000000000000 ;
        1814:  q   <=  32'b00000000000000000000000000000000 ;
        1815:  q   <=  32'b00000000000000000000000000000000 ;
        1816:  q   <=  32'b00000000000000000000000000000000 ;
        1817:  q   <=  32'b00000000000000000000000000000000 ;
        1818:  q   <=  32'b00000000000000000000000000000000 ;
        1819:  q   <=  32'b00000000000000000000000000000000 ;
        1820:  q   <=  32'b00000000000000000000000000000000 ;
        1821:  q   <=  32'b00000000000000000000000000000000 ;
        1822:  q   <=  32'b00000000000000000000000000000000 ;
        1823:  q   <=  32'b00000000000000000000000000000000 ;
        1824:  q   <=  32'b00000000000000000000000000000000 ;
        1825:  q   <=  32'b00000000000000000000000000000000 ;
        1826:  q   <=  32'b00000000000000000000000000000000 ;
        1827:  q   <=  32'b00000000000000000000000000000000 ;
        1828:  q   <=  32'b00000000000000000000000000000000 ;
        1829:  q   <=  32'b00000000000000000000000000000000 ;
        1830:  q   <=  32'b00000000000000000000000000000000 ;
        1831:  q   <=  32'b00000000000000000000000000000000 ;
        1832:  q   <=  32'b00000000000000000000000000000000 ;
        1833:  q   <=  32'b00000000000000000000000000000000 ;
        1834:  q   <=  32'b00000000000000000000000000000000 ;
        1835:  q   <=  32'b00000000000000000000000000000000 ;
        1836:  q   <=  32'b00000000000000000000000000000000 ;
        1837:  q   <=  32'b00000000000000000000000000000000 ;
        1838:  q   <=  32'b00000000000000000000000000000000 ;
        1839:  q   <=  32'b00000000000000000000000000000000 ;
        1840:  q   <=  32'b00000000000000000000000000000000 ;
        1841:  q   <=  32'b00000000000000000000000000000000 ;
        1842:  q   <=  32'b00000000000000000000000000000000 ;
        1843:  q   <=  32'b00000000000000000000000000000000 ;
        1844:  q   <=  32'b00000000000000000000000000000000 ;
        1845:  q   <=  32'b00000000000000000000000000000000 ;
        1846:  q   <=  32'b00000000000000000000000000000000 ;
        1847:  q   <=  32'b00000000000000000000000000000000 ;
        1848:  q   <=  32'b00000000000000000000000000000000 ;
        1849:  q   <=  32'b00000000000000000000000000000000 ;
        1850:  q   <=  32'b00000000000000000000000000000000 ;
        1851:  q   <=  32'b00000000000000000000000000000000 ;
        1852:  q   <=  32'b00000000000000000000000000000000 ;
        1853:  q   <=  32'b00000000000000000000000000000000 ;
        1854:  q   <=  32'b00000000000000000000000000000000 ;
        1855:  q   <=  32'b00000000000000000000000000000000 ;
        1856:  q   <=  32'b00000000000000000000000000000000 ;
        1857:  q   <=  32'b00000000000000000000000000000000 ;
        1858:  q   <=  32'b00000000000000000000000000000000 ;
        1859:  q   <=  32'b00000000000000000000000000000000 ;
        1860:  q   <=  32'b00000000000000000000000000000000 ;
        1861:  q   <=  32'b00000000000000000000000000000000 ;
        1862:  q   <=  32'b00000000000000000000000000000000 ;
        1863:  q   <=  32'b00000000000000000000000000000000 ;
        1864:  q   <=  32'b00000000000000000000000000000000 ;
        1865:  q   <=  32'b00000000000000000000000000000000 ;
        1866:  q   <=  32'b00000000000000000000000000000000 ;
        1867:  q   <=  32'b00000000000000000000000000000000 ;
        1868:  q   <=  32'b00000000000000000000000000000000 ;
        1869:  q   <=  32'b00000000000000000000000000000000 ;
        1870:  q   <=  32'b00000000000000000000000000000000 ;
        1871:  q   <=  32'b00000000000000000000000000000000 ;
        1872:  q   <=  32'b00000000000000000000000000000000 ;
        1873:  q   <=  32'b00000000000000000000000000000000 ;
        1874:  q   <=  32'b00000000000000000000000000000000 ;
        1875:  q   <=  32'b00000000000000000000000000000000 ;
        1876:  q   <=  32'b00000000000000000000000000000000 ;
        1877:  q   <=  32'b00000000000000000000000000000000 ;
        1878:  q   <=  32'b00000000000000000000000000000000 ;
        1879:  q   <=  32'b00000000000000000000000000000000 ;
        1880:  q   <=  32'b00000000000000000000000000000000 ;
        1881:  q   <=  32'b00000000000000000000000000000000 ;
        1882:  q   <=  32'b00000000000000000000000000000000 ;
        1883:  q   <=  32'b00000000000000000000000000000000 ;
        1884:  q   <=  32'b00000000000000000000000000000000 ;
        1885:  q   <=  32'b00000000000000000000000000000000 ;
        1886:  q   <=  32'b00000000000000000000000000000000 ;
        1887:  q   <=  32'b00000000000000000000000000000000 ;
        1888:  q   <=  32'b00000000000000000000000000000000 ;
        1889:  q   <=  32'b00000000000000000000000000000000 ;
        1890:  q   <=  32'b00000000000000000000000000000000 ;
        1891:  q   <=  32'b00000000000000000000000000000000 ;
        1892:  q   <=  32'b00000000000000000000000000000000 ;
        1893:  q   <=  32'b00000000000000000000000000000000 ;
        1894:  q   <=  32'b00000000000000000000000000000000 ;
        1895:  q   <=  32'b00000000000000000000000000000000 ;
        1896:  q   <=  32'b00000000000000000000000000000000 ;
        1897:  q   <=  32'b00000000000000000000000000000000 ;
        1898:  q   <=  32'b00000000000000000000000000000000 ;
        1899:  q   <=  32'b00000000000000000000000000000000 ;
        1900:  q   <=  32'b00000000000000000000000000000000 ;
        1901:  q   <=  32'b00000000000000000000000000000000 ;
        1902:  q   <=  32'b00000000000000000000000000000000 ;
        1903:  q   <=  32'b00000000000000000000000000000000 ;
        1904:  q   <=  32'b00000000000000000000000000000000 ;
        1905:  q   <=  32'b00000000000000000000000000000000 ;
        1906:  q   <=  32'b00000000000000000000000000000000 ;
        1907:  q   <=  32'b00000000000000000000000000000000 ;
        1908:  q   <=  32'b00000000000000000000000000000000 ;
        1909:  q   <=  32'b00000000000000000000000000000000 ;
        1910:  q   <=  32'b00000000000000000000000000000000 ;
        1911:  q   <=  32'b00000000000000000000000000000000 ;
        1912:  q   <=  32'b00000000000000000000000000000000 ;
        1913:  q   <=  32'b00000000000000000000000000000000 ;
        1914:  q   <=  32'b00000000000000000000000000000000 ;
        1915:  q   <=  32'b00000000000000000000000000000000 ;
        1916:  q   <=  32'b00000000000000000000000000000000 ;
        1917:  q   <=  32'b00000000000000000000000000000000 ;
        1918:  q   <=  32'b00000000000000000000000000000000 ;
        1919:  q   <=  32'b00000000000000000000000000000000 ;
        1920:  q   <=  32'b00000000000000000000000000000000 ;
        1921:  q   <=  32'b00000000000000000000000000000000 ;
        1922:  q   <=  32'b00000000000000000000000000000000 ;
        1923:  q   <=  32'b00000000000000000000000000000000 ;
        1924:  q   <=  32'b00000000000000000000000000000000 ;
        1925:  q   <=  32'b00000000000000000000000000000000 ;
        1926:  q   <=  32'b00000000000000000000000000000000 ;
        1927:  q   <=  32'b00000000000000000000000000000000 ;
        1928:  q   <=  32'b00000000000000000000000000000000 ;
        1929:  q   <=  32'b00000000000000000000000000000000 ;
        1930:  q   <=  32'b00000000000000000000000000000000 ;
        1931:  q   <=  32'b00000000000000000000000000000000 ;
        1932:  q   <=  32'b00000000000000000000000000000000 ;
        1933:  q   <=  32'b00000000000000000000000000000000 ;
        1934:  q   <=  32'b00000000000000000000000000000000 ;
        1935:  q   <=  32'b00000000000000000000000000000000 ;
        1936:  q   <=  32'b00000000000000000000000000000000 ;
        1937:  q   <=  32'b00000000000000000000000000000000 ;
        1938:  q   <=  32'b00000000000000000000000000000000 ;
        1939:  q   <=  32'b00000000000000000000000000000000 ;
        1940:  q   <=  32'b00000000000000000000000000000000 ;
        1941:  q   <=  32'b00000000000000000000000000000000 ;
        1942:  q   <=  32'b00000000000000000000000000000000 ;
        1943:  q   <=  32'b00000000000000000000000000000000 ;
        1944:  q   <=  32'b00000000000000000000000000000000 ;
        1945:  q   <=  32'b00000000000000000000000000000000 ;
        1946:  q   <=  32'b00000000000000000000000000000000 ;
        1947:  q   <=  32'b00000000000000000000000000000000 ;
        1948:  q   <=  32'b00000000000000000000000000000000 ;
        1949:  q   <=  32'b00000000000000000000000000000000 ;
        1950:  q   <=  32'b00000000000000000000000000000000 ;
        1951:  q   <=  32'b00000000000000000000000000000000 ;
        1952:  q   <=  32'b00000000000000000000000000000000 ;
        1953:  q   <=  32'b00000000000000000000000000000000 ;
        1954:  q   <=  32'b00000000000000000000000000000000 ;
        1955:  q   <=  32'b00000000000000000000000000000000 ;
        1956:  q   <=  32'b00000000000000000000000000000000 ;
        1957:  q   <=  32'b00000000000000000000000000000000 ;
        1958:  q   <=  32'b00000000000000000000000000000000 ;
        1959:  q   <=  32'b00000000000000000000000000000000 ;
        1960:  q   <=  32'b00000000000000000000000000000000 ;
        1961:  q   <=  32'b00000000000000000000000000000000 ;
        1962:  q   <=  32'b00000000000000000000000000000000 ;
        1963:  q   <=  32'b00000000000000000000000000000000 ;
        1964:  q   <=  32'b00000000000000000000000000000000 ;
        1965:  q   <=  32'b00111100111000000011011111000110 ;
        1966:  q   <=  32'b00111110100110110011110111000111 ;
        1967:  q   <=  32'b00111111000100111100001110110010 ;
        1968:  q   <=  32'b00111111010110010111000101011110 ;
        1969:  q   <=  32'b00111111100011110101010010001001 ;
        1970:  q   <=  32'b00111111101100011011010111111111 ;
        1971:  q   <=  32'b00111111110100111101110110100010 ;
        1972:  q   <=  32'b00111111111101011100110000000101 ;
        1973:  q   <=  32'b00111111111010000111111001001000 ;
        1974:  q   <=  32'b00111111110001110000000010111010 ;
        1975:  q   <=  32'b00111111101001011011101011000100 ;
        1976:  q   <=  32'b00111111100001001010101111011100 ;
        1977:  q   <=  32'b00111111010001111010011011110011 ;
        1978:  q   <=  32'b00111111000001100110001000101100 ;
        1979:  q   <=  32'b00111110100010110001000010110101 ;
        1980:  q   <=  32'b00111100101000110000111011110110 ;
        1981:  q   <=  32'b00000000000000000000000000000000 ;
        1982:  q   <=  32'b00000000000000000000000000000000 ;
        1983:  q   <=  32'b00000000000000000000000000000000 ;
        1984:  q   <=  32'b00000000000000000000000000000000 ;
        1985:  q   <=  32'b00000000000000000000000000000000 ;
        1986:  q   <=  32'b00000000000000000000000000000000 ;
        1987:  q   <=  32'b00000000000000000000000000000000 ;
        1988:  q   <=  32'b00000000000000000000000000000000 ;
        1989:  q   <=  32'b00000000000000000000000000000000 ;
        1990:  q   <=  32'b00000000000000000000000000000000 ;
        1991:  q   <=  32'b00000000000000000000000000000000 ;
        1992:  q   <=  32'b00000000000000000000000000000000 ;
        1993:  q   <=  32'b00000000000000000000000000000000 ;
        1994:  q   <=  32'b00000000000000000000000000000000 ;
        1995:  q   <=  32'b00000000000000000000000000000000 ;
        1996:  q   <=  32'b00000000000000000000000000000000 ;
        1997:  q   <=  32'b00000000000000000000000000000000 ;
        1998:  q   <=  32'b00000000000000000000000000000000 ;
        1999:  q   <=  32'b00000000000000000000000000000000 ;
        2000:  q   <=  32'b00000000000000000000000000000000 ;
        2001:  q   <=  32'b00000000000000000000000000000000 ;
        2002:  q   <=  32'b00000000000000000000000000000000 ;
        2003:  q   <=  32'b00000000000000000000000000000000 ;
        2004:  q   <=  32'b00000000000000000000000000000000 ;
        2005:  q   <=  32'b00000000000000000000000000000000 ;
        2006:  q   <=  32'b00000000000000000000000000000000 ;
        2007:  q   <=  32'b00000000000000000000000000000000 ;
        2008:  q   <=  32'b00000000000000000000000000000000 ;
        2009:  q   <=  32'b00000000000000000000000000000000 ;
        2010:  q   <=  32'b00000000000000000000000000000000 ;
        2011:  q   <=  32'b00000000000000000000000000000000 ;
        2012:  q   <=  32'b00000000000000000000000000000000 ;
        2013:  q   <=  32'b00000000000000000000000000000000 ;
        2014:  q   <=  32'b00000000000000000000000000000000 ;
        2015:  q   <=  32'b00000000000000000000000000000000 ;
        2016:  q   <=  32'b00000000000000000000000000000000 ;
        2017:  q   <=  32'b00000000000000000000000000000000 ;
        2018:  q   <=  32'b00000000000000000000000000000000 ;
        2019:  q   <=  32'b00000000000000000000000000000000 ;
        2020:  q   <=  32'b00000000000000000000000000000000 ;
        2021:  q   <=  32'b00000000000000000000000000000000 ;
        2022:  q   <=  32'b00000000000000000000000000000000 ;
        2023:  q   <=  32'b00000000000000000000000000000000 ;
        2024:  q   <=  32'b00000000000000000000000000000000 ;
        2025:  q   <=  32'b00000000000000000000000000000000 ;
        2026:  q   <=  32'b00000000000000000000000000000000 ;
        2027:  q   <=  32'b00000000000000000000000000000000 ;
        2028:  q   <=  32'b00000000000000000000000000000000 ;
        2029:  q   <=  32'b00000000000000000000000000000000 ;
        2030:  q   <=  32'b00000000000000000000000000000000 ;
        2031:  q   <=  32'b00000000000000000000000000000000 ;
        2032:  q   <=  32'b00000000000000000000000000000000 ;
        2033:  q   <=  32'b00000000000000000000000000000000 ;
        2034:  q   <=  32'b00000000000000000000000000000000 ;
        2035:  q   <=  32'b00000000000000000000000000000000 ;
        2036:  q   <=  32'b00000000000000000000000000000000 ;
        2037:  q   <=  32'b00000000000000000000000000000000 ;
        2038:  q   <=  32'b00000000000000000000000000000000 ;
        2039:  q   <=  32'b00000000000000000000000000000000 ;
        2040:  q   <=  32'b00000000000000000000000000000000 ;
        2041:  q   <=  32'b00000000000000000000000000000000 ;
        2042:  q   <=  32'b00000000000000000000000000000000 ;
        2043:  q   <=  32'b00000000000000000000000000000000 ;
        2044:  q   <=  32'b00000000000000000000000000000000 ;
        2045:  q   <=  32'b00000000000000000000000000000000 ;
        2046:  q   <=  32'b00000000000000000000000000000000 ;
        2047:  q   <=  32'b00000000000000000000000000000000 ;
        2048:  q   <=  32'b00000000000000000000000000000000 ;
        2049:  q   <=  32'b00000000000000000000000000000000 ;
        2050:  q   <=  32'b00000000000000000000000000000000 ;
        2051:  q   <=  32'b00000000000000000000000000000000 ;
        2052:  q   <=  32'b00000000000000000000000000000000 ;
        2053:  q   <=  32'b00000000000000000000000000000000 ;
        2054:  q   <=  32'b00000000000000000000000000000000 ;
        2055:  q   <=  32'b00000000000000000000000000000000 ;
        2056:  q   <=  32'b00000000000000000000000000000000 ;
        2057:  q   <=  32'b00000000000000000000000000000000 ;
        2058:  q   <=  32'b00000000000000000000000000000000 ;
        2059:  q   <=  32'b00000000000000000000000000000000 ;
        2060:  q   <=  32'b00000000000000000000000000000000 ;
        2061:  q   <=  32'b00000000000000000000000000000000 ;
        2062:  q   <=  32'b00000000000000000000000000000000 ;
        2063:  q   <=  32'b00000000000000000000000000000000 ;
        2064:  q   <=  32'b00000000000000000000000000000000 ;
        2065:  q   <=  32'b00000000000000000000000000000000 ;
        2066:  q   <=  32'b00000000000000000000000000000000 ;
        2067:  q   <=  32'b00000000000000000000000000000000 ;
        2068:  q   <=  32'b00000000000000000000000000000000 ;
        2069:  q   <=  32'b00000000000000000000000000000000 ;
        2070:  q   <=  32'b00000000000000000000000000000000 ;
        2071:  q   <=  32'b00000000000000000000000000000000 ;
        2072:  q   <=  32'b00000000000000000000000000000000 ;
        2073:  q   <=  32'b00000000000000000000000000000000 ;
        2074:  q   <=  32'b00000000000000000000000000000000 ;
        2075:  q   <=  32'b00000000000000000000000000000000 ;
        2076:  q   <=  32'b00000000000000000000000000000000 ;
        2077:  q   <=  32'b00000000000000000000000000000000 ;
        2078:  q   <=  32'b00000000000000000000000000000000 ;
        2079:  q   <=  32'b00000000000000000000000000000000 ;
        2080:  q   <=  32'b00000000000000000000000000000000 ;
        2081:  q   <=  32'b00000000000000000000000000000000 ;
        2082:  q   <=  32'b00000000000000000000000000000000 ;
        2083:  q   <=  32'b00000000000000000000000000000000 ;
        2084:  q   <=  32'b00000000000000000000000000000000 ;
        2085:  q   <=  32'b00000000000000000000000000000000 ;
        2086:  q   <=  32'b00000000000000000000000000000000 ;
        2087:  q   <=  32'b00000000000000000000000000000000 ;
        2088:  q   <=  32'b00000000000000000000000000000000 ;
        2089:  q   <=  32'b00000000000000000000000000000000 ;
        2090:  q   <=  32'b00000000000000000000000000000000 ;
        2091:  q   <=  32'b00000000000000000000000000000000 ;
        2092:  q   <=  32'b00000000000000000000000000000000 ;
        2093:  q   <=  32'b00000000000000000000000000000000 ;
        2094:  q   <=  32'b00000000000000000000000000000000 ;
        2095:  q   <=  32'b00000000000000000000000000000000 ;
        2096:  q   <=  32'b00000000000000000000000000000000 ;
        2097:  q   <=  32'b00000000000000000000000000000000 ;
        2098:  q   <=  32'b00000000000000000000000000000000 ;
        2099:  q   <=  32'b00000000000000000000000000000000 ;
        2100:  q   <=  32'b00000000000000000000000000000000 ;
        2101:  q   <=  32'b00000000000000000000000000000000 ;
        2102:  q   <=  32'b00000000000000000000000000000000 ;
        2103:  q   <=  32'b00000000000000000000000000000000 ;
        2104:  q   <=  32'b00000000000000000000000000000000 ;
        2105:  q   <=  32'b00000000000000000000000000000000 ;
        2106:  q   <=  32'b00000000000000000000000000000000 ;
        2107:  q   <=  32'b00000000000000000000000000000000 ;
        2108:  q   <=  32'b00000000000000000000000000000000 ;
        2109:  q   <=  32'b00000000000000000000000000000000 ;
        2110:  q   <=  32'b00000000000000000000000000000000 ;
        2111:  q   <=  32'b00000000000000000000000000000000 ;
        2112:  q   <=  32'b00000000000000000000000000000000 ;
        2113:  q   <=  32'b00000000000000000000000000000000 ;
        2114:  q   <=  32'b00000000000000000000000000000000 ;
        2115:  q   <=  32'b00000000000000000000000000000000 ;
        2116:  q   <=  32'b00000000000000000000000000000000 ;
        2117:  q   <=  32'b00000000000000000000000000000000 ;
        2118:  q   <=  32'b00000000000000000000000000000000 ;
        2119:  q   <=  32'b00000000000000000000000000000000 ;
        2120:  q   <=  32'b00000000000000000000000000000000 ;
        2121:  q   <=  32'b00000000000000000000000000000000 ;
        2122:  q   <=  32'b00000000000000000000000000000000 ;
        2123:  q   <=  32'b00000000000000000000000000000000 ;
        2124:  q   <=  32'b00000000000000000000000000000000 ;
        2125:  q   <=  32'b00000000000000000000000000000000 ;
        2126:  q   <=  32'b00000000000000000000000000000000 ;
        2127:  q   <=  32'b00000000000000000000000000000000 ;
        2128:  q   <=  32'b00000000000000000000000000000000 ;
        2129:  q   <=  32'b00000000000000000000000000000000 ;
        2130:  q   <=  32'b00000000000000000000000000000000 ;
        2131:  q   <=  32'b00000000000000000000000000000000 ;
        2132:  q   <=  32'b00000000000000000000000000000000 ;
        2133:  q   <=  32'b00000000000000000000000000000000 ;
        2134:  q   <=  32'b00000000000000000000000000000000 ;
        2135:  q   <=  32'b00000000000000000000000000000000 ;
        2136:  q   <=  32'b00000000000000000000000000000000 ;
        2137:  q   <=  32'b00000000000000000000000000000000 ;
        2138:  q   <=  32'b00000000000000000000000000000000 ;
        2139:  q   <=  32'b00000000000000000000000000000000 ;
        2140:  q   <=  32'b00000000000000000000000000000000 ;
        2141:  q   <=  32'b00000000000000000000000000000000 ;
        2142:  q   <=  32'b00000000000000000000000000000000 ;
        2143:  q   <=  32'b00000000000000000000000000000000 ;
        2144:  q   <=  32'b00000000000000000000000000000000 ;
        2145:  q   <=  32'b00000000000000000000000000000000 ;
        2146:  q   <=  32'b00000000000000000000000000000000 ;
        2147:  q   <=  32'b00000000000000000000000000000000 ;
        2148:  q   <=  32'b00000000000000000000000000000000 ;
        2149:  q   <=  32'b00000000000000000000000000000000 ;
        2150:  q   <=  32'b00000000000000000000000000000000 ;
        2151:  q   <=  32'b00000000000000000000000000000000 ;
        2152:  q   <=  32'b00000000000000000000000000000000 ;
        2153:  q   <=  32'b00000000000000000000000000000000 ;
        2154:  q   <=  32'b00000000000000000000000000000000 ;
        2155:  q   <=  32'b00000000000000000000000000000000 ;
        2156:  q   <=  32'b00000000000000000000000000000000 ;
        2157:  q   <=  32'b00000000000000000000000000000000 ;
        2158:  q   <=  32'b00000000000000000000000000000000 ;
        2159:  q   <=  32'b00000000000000000000000000000000 ;
        2160:  q   <=  32'b00000000000000000000000000000000 ;
        2161:  q   <=  32'b00000000000000000000000000000000 ;
        2162:  q   <=  32'b00000000000000000000000000000000 ;
        2163:  q   <=  32'b00000000000000000000000000000000 ;
        2164:  q   <=  32'b00000000000000000000000000000000 ;
        2165:  q   <=  32'b00000000000000000000000000000000 ;
        2166:  q   <=  32'b00000000000000000000000000000000 ;
        2167:  q   <=  32'b00000000000000000000000000000000 ;
        2168:  q   <=  32'b00000000000000000000000000000000 ;
        2169:  q   <=  32'b00000000000000000000000000000000 ;
        2170:  q   <=  32'b00000000000000000000000000000000 ;
        2171:  q   <=  32'b00000000000000000000000000000000 ;
        2172:  q   <=  32'b00000000000000000000000000000000 ;
        2173:  q   <=  32'b00000000000000000000000000000000 ;
        2174:  q   <=  32'b00000000000000000000000000000000 ;
        2175:  q   <=  32'b00000000000000000000000000000000 ;
        2176:  q   <=  32'b00000000000000000000000000000000 ;
        2177:  q   <=  32'b00000000000000000000000000000000 ;
        2178:  q   <=  32'b00000000000000000000000000000000 ;
        2179:  q   <=  32'b00000000000000000000000000000000 ;
        2180:  q   <=  32'b00000000000000000000000000000000 ;
        2181:  q   <=  32'b00000000000000000000000000000000 ;
        2182:  q   <=  32'b00000000000000000000000000000000 ;
        2183:  q   <=  32'b00000000000000000000000000000000 ;
        2184:  q   <=  32'b00000000000000000000000000000000 ;
        2185:  q   <=  32'b00000000000000000000000000000000 ;
        2186:  q   <=  32'b00000000000000000000000000000000 ;
        2187:  q   <=  32'b00000000000000000000000000000000 ;
        2188:  q   <=  32'b00000000000000000000000000000000 ;
        2189:  q   <=  32'b00000000000000000000000000000000 ;
        2190:  q   <=  32'b00000000000000000000000000000000 ;
        2191:  q   <=  32'b00000000000000000000000000000000 ;
        2192:  q   <=  32'b00000000000000000000000000000000 ;
        2193:  q   <=  32'b00000000000000000000000000000000 ;
        2194:  q   <=  32'b00000000000000000000000000000000 ;
        2195:  q   <=  32'b00000000000000000000000000000000 ;
        2196:  q   <=  32'b00000000000000000000000000000000 ;
        2197:  q   <=  32'b00000000000000000000000000000000 ;
        2198:  q   <=  32'b00000000000000000000000000000000 ;
        2199:  q   <=  32'b00000000000000000000000000000000 ;
        2200:  q   <=  32'b00000000000000000000000000000000 ;
        2201:  q   <=  32'b00000000000000000000000000000000 ;
        2202:  q   <=  32'b00000000000000000000000000000000 ;
        2203:  q   <=  32'b00000000000000000000000000000000 ;
        2204:  q   <=  32'b00000000000000000000000000000000 ;
        2205:  q   <=  32'b00000000000000000000000000000000 ;
        2206:  q   <=  32'b00000000000000000000000000000000 ;
        2207:  q   <=  32'b00000000000000000000000000000000 ;
        2208:  q   <=  32'b00000000000000000000000000000000 ;
        2209:  q   <=  32'b00000000000000000000000000000000 ;
        2210:  q   <=  32'b00000000000000000000000000000000 ;
        2211:  q   <=  32'b00000000000000000000000000000000 ;
        2212:  q   <=  32'b00000000000000000000000000000000 ;
        2213:  q   <=  32'b00000000000000000000000000000000 ;
        2214:  q   <=  32'b00000000000000000000000000000000 ;
        2215:  q   <=  32'b00000000000000000000000000000000 ;
        2216:  q   <=  32'b00000000000000000000000000000000 ;
        2217:  q   <=  32'b00000000000000000000000000000000 ;
        2218:  q   <=  32'b00000000000000000000000000000000 ;
        2219:  q   <=  32'b00000000000000000000000000000000 ;
        2220:  q   <=  32'b00000000000000000000000000000000 ;
        2221:  q   <=  32'b00000000000000000000000000000000 ;
        2222:  q   <=  32'b00000000000000000000000000000000 ;
        2223:  q   <=  32'b00000000000000000000000000000000 ;
        2224:  q   <=  32'b00000000000000000000000000000000 ;
        2225:  q   <=  32'b00000000000000000000000000000000 ;
        2226:  q   <=  32'b00000000000000000000000000000000 ;
        2227:  q   <=  32'b00000000000000000000000000000000 ;
        2228:  q   <=  32'b00000000000000000000000000000000 ;
        2229:  q   <=  32'b00111110001111000000110110111001 ;
        2230:  q   <=  32'b00111110111000111111110100010100 ;
        2231:  q   <=  32'b00111111001101001000101001110110 ;
        2232:  q   <=  32'b00111111011101101010100001000110 ;
        2233:  q   <=  32'b00111111100111000010110010000110 ;
        2234:  q   <=  32'b00111111101111001100111011101001 ;
        2235:  q   <=  32'b00111111110111010011101111010010 ;
        2236:  q   <=  32'b00111111111111010111001111000100 ;
        2237:  q   <=  32'b00111111111000101000100011000000 ;
        2238:  q   <=  32'b00111111110000101011100100111011 ;
        2239:  q   <=  32'b00111111101000110001110100101110 ;
        2240:  q   <=  32'b00111111100000111011010000011100 ;
        2241:  q   <=  32'b00111111010010001111101100011000 ;
        2242:  q   <=  32'b00111111000010101111001000000110 ;
        2243:  q   <=  32'b00111110100110101001100000100101 ;
        2244:  q   <=  32'b00111101100000000100001010001000 ;
        2245:  q   <=  32'b00000000000000000000000000000000 ;
        2246:  q   <=  32'b00000000000000000000000000000000 ;
        2247:  q   <=  32'b00000000000000000000000000000000 ;
        2248:  q   <=  32'b00000000000000000000000000000000 ;
        2249:  q   <=  32'b00000000000000000000000000000000 ;
        2250:  q   <=  32'b00000000000000000000000000000000 ;
        2251:  q   <=  32'b00000000000000000000000000000000 ;
        2252:  q   <=  32'b00000000000000000000000000000000 ;
        2253:  q   <=  32'b00000000000000000000000000000000 ;
        2254:  q   <=  32'b00000000000000000000000000000000 ;
        2255:  q   <=  32'b00000000000000000000000000000000 ;
        2256:  q   <=  32'b00000000000000000000000000000000 ;
        2257:  q   <=  32'b00000000000000000000000000000000 ;
        2258:  q   <=  32'b00000000000000000000000000000000 ;
        2259:  q   <=  32'b00000000000000000000000000000000 ;
        2260:  q   <=  32'b00000000000000000000000000000000 ;
        2261:  q   <=  32'b00000000000000000000000000000000 ;
        2262:  q   <=  32'b00000000000000000000000000000000 ;
        2263:  q   <=  32'b00000000000000000000000000000000 ;
        2264:  q   <=  32'b00000000000000000000000000000000 ;
        2265:  q   <=  32'b00000000000000000000000000000000 ;
        2266:  q   <=  32'b00000000000000000000000000000000 ;
        2267:  q   <=  32'b00000000000000000000000000000000 ;
        2268:  q   <=  32'b00000000000000000000000000000000 ;
        2269:  q   <=  32'b00000000000000000000000000000000 ;
        2270:  q   <=  32'b00000000000000000000000000000000 ;
        2271:  q   <=  32'b00000000000000000000000000000000 ;
        2272:  q   <=  32'b00000000000000000000000000000000 ;
        2273:  q   <=  32'b00000000000000000000000000000000 ;
        2274:  q   <=  32'b00000000000000000000000000000000 ;
        2275:  q   <=  32'b00000000000000000000000000000000 ;
        2276:  q   <=  32'b00000000000000000000000000000000 ;
        2277:  q   <=  32'b00000000000000000000000000000000 ;
        2278:  q   <=  32'b00000000000000000000000000000000 ;
        2279:  q   <=  32'b00000000000000000000000000000000 ;
        2280:  q   <=  32'b00000000000000000000000000000000 ;
        2281:  q   <=  32'b00000000000000000000000000000000 ;
        2282:  q   <=  32'b00000000000000000000000000000000 ;
        2283:  q   <=  32'b00000000000000000000000000000000 ;
        2284:  q   <=  32'b00000000000000000000000000000000 ;
        2285:  q   <=  32'b00000000000000000000000000000000 ;
        2286:  q   <=  32'b00000000000000000000000000000000 ;
        2287:  q   <=  32'b00000000000000000000000000000000 ;
        2288:  q   <=  32'b00000000000000000000000000000000 ;
        2289:  q   <=  32'b00000000000000000000000000000000 ;
        2290:  q   <=  32'b00000000000000000000000000000000 ;
        2291:  q   <=  32'b00000000000000000000000000000000 ;
        2292:  q   <=  32'b00000000000000000000000000000000 ;
        2293:  q   <=  32'b00000000000000000000000000000000 ;
        2294:  q   <=  32'b00000000000000000000000000000000 ;
        2295:  q   <=  32'b00000000000000000000000000000000 ;
        2296:  q   <=  32'b00000000000000000000000000000000 ;
        2297:  q   <=  32'b00000000000000000000000000000000 ;
        2298:  q   <=  32'b00000000000000000000000000000000 ;
        2299:  q   <=  32'b00000000000000000000000000000000 ;
        2300:  q   <=  32'b00000000000000000000000000000000 ;
        2301:  q   <=  32'b00000000000000000000000000000000 ;
        2302:  q   <=  32'b00000000000000000000000000000000 ;
        2303:  q   <=  32'b00000000000000000000000000000000 ;
        2304:  q   <=  32'b00000000000000000000000000000000 ;
        2305:  q   <=  32'b00000000000000000000000000000000 ;
        2306:  q   <=  32'b00000000000000000000000000000000 ;
        2307:  q   <=  32'b00000000000000000000000000000000 ;
        2308:  q   <=  32'b00000000000000000000000000000000 ;
        2309:  q   <=  32'b00000000000000000000000000000000 ;
        2310:  q   <=  32'b00000000000000000000000000000000 ;
        2311:  q   <=  32'b00000000000000000000000000000000 ;
        2312:  q   <=  32'b00000000000000000000000000000000 ;
        2313:  q   <=  32'b00000000000000000000000000000000 ;
        2314:  q   <=  32'b00000000000000000000000000000000 ;
        2315:  q   <=  32'b00000000000000000000000000000000 ;
        2316:  q   <=  32'b00000000000000000000000000000000 ;
        2317:  q   <=  32'b00000000000000000000000000000000 ;
        2318:  q   <=  32'b00000000000000000000000000000000 ;
        2319:  q   <=  32'b00000000000000000000000000000000 ;
        2320:  q   <=  32'b00000000000000000000000000000000 ;
        2321:  q   <=  32'b00000000000000000000000000000000 ;
        2322:  q   <=  32'b00000000000000000000000000000000 ;
        2323:  q   <=  32'b00000000000000000000000000000000 ;
        2324:  q   <=  32'b00000000000000000000000000000000 ;
        2325:  q   <=  32'b00000000000000000000000000000000 ;
        2326:  q   <=  32'b00000000000000000000000000000000 ;
        2327:  q   <=  32'b00000000000000000000000000000000 ;
        2328:  q   <=  32'b00000000000000000000000000000000 ;
        2329:  q   <=  32'b00000000000000000000000000000000 ;
        2330:  q   <=  32'b00000000000000000000000000000000 ;
        2331:  q   <=  32'b00000000000000000000000000000000 ;
        2332:  q   <=  32'b00000000000000000000000000000000 ;
        2333:  q   <=  32'b00000000000000000000000000000000 ;
        2334:  q   <=  32'b00000000000000000000000000000000 ;
        2335:  q   <=  32'b00000000000000000000000000000000 ;
        2336:  q   <=  32'b00000000000000000000000000000000 ;
        2337:  q   <=  32'b00000000000000000000000000000000 ;
        2338:  q   <=  32'b00000000000000000000000000000000 ;
        2339:  q   <=  32'b00000000000000000000000000000000 ;
        2340:  q   <=  32'b00000000000000000000000000000000 ;
        2341:  q   <=  32'b00000000000000000000000000000000 ;
        2342:  q   <=  32'b00000000000000000000000000000000 ;
        2343:  q   <=  32'b00000000000000000000000000000000 ;
        2344:  q   <=  32'b00000000000000000000000000000000 ;
        2345:  q   <=  32'b00000000000000000000000000000000 ;
        2346:  q   <=  32'b00000000000000000000000000000000 ;
        2347:  q   <=  32'b00000000000000000000000000000000 ;
        2348:  q   <=  32'b00000000000000000000000000000000 ;
        2349:  q   <=  32'b00000000000000000000000000000000 ;
        2350:  q   <=  32'b00000000000000000000000000000000 ;
        2351:  q   <=  32'b00000000000000000000000000000000 ;
        2352:  q   <=  32'b00000000000000000000000000000000 ;
        2353:  q   <=  32'b00000000000000000000000000000000 ;
        2354:  q   <=  32'b00000000000000000000000000000000 ;
        2355:  q   <=  32'b00000000000000000000000000000000 ;
        2356:  q   <=  32'b00000000000000000000000000000000 ;
        2357:  q   <=  32'b00000000000000000000000000000000 ;
        2358:  q   <=  32'b00000000000000000000000000000000 ;
        2359:  q   <=  32'b00000000000000000000000000000000 ;
        2360:  q   <=  32'b00000000000000000000000000000000 ;
        2361:  q   <=  32'b00000000000000000000000000000000 ;
        2362:  q   <=  32'b00000000000000000000000000000000 ;
        2363:  q   <=  32'b00000000000000000000000000000000 ;
        2364:  q   <=  32'b00000000000000000000000000000000 ;
        2365:  q   <=  32'b00000000000000000000000000000000 ;
        2366:  q   <=  32'b00000000000000000000000000000000 ;
        2367:  q   <=  32'b00000000000000000000000000000000 ;
        2368:  q   <=  32'b00000000000000000000000000000000 ;
        2369:  q   <=  32'b00000000000000000000000000000000 ;
        2370:  q   <=  32'b00000000000000000000000000000000 ;
        2371:  q   <=  32'b00000000000000000000000000000000 ;
        2372:  q   <=  32'b00000000000000000000000000000000 ;
        2373:  q   <=  32'b00000000000000000000000000000000 ;
        2374:  q   <=  32'b00000000000000000000000000000000 ;
        2375:  q   <=  32'b00000000000000000000000000000000 ;
        2376:  q   <=  32'b00000000000000000000000000000000 ;
        2377:  q   <=  32'b00000000000000000000000000000000 ;
        2378:  q   <=  32'b00000000000000000000000000000000 ;
        2379:  q   <=  32'b00000000000000000000000000000000 ;
        2380:  q   <=  32'b00000000000000000000000000000000 ;
        2381:  q   <=  32'b00000000000000000000000000000000 ;
        2382:  q   <=  32'b00000000000000000000000000000000 ;
        2383:  q   <=  32'b00000000000000000000000000000000 ;
        2384:  q   <=  32'b00000000000000000000000000000000 ;
        2385:  q   <=  32'b00000000000000000000000000000000 ;
        2386:  q   <=  32'b00000000000000000000000000000000 ;
        2387:  q   <=  32'b00000000000000000000000000000000 ;
        2388:  q   <=  32'b00000000000000000000000000000000 ;
        2389:  q   <=  32'b00000000000000000000000000000000 ;
        2390:  q   <=  32'b00000000000000000000000000000000 ;
        2391:  q   <=  32'b00000000000000000000000000000000 ;
        2392:  q   <=  32'b00000000000000000000000000000000 ;
        2393:  q   <=  32'b00000000000000000000000000000000 ;
        2394:  q   <=  32'b00000000000000000000000000000000 ;
        2395:  q   <=  32'b00000000000000000000000000000000 ;
        2396:  q   <=  32'b00000000000000000000000000000000 ;
        2397:  q   <=  32'b00000000000000000000000000000000 ;
        2398:  q   <=  32'b00000000000000000000000000000000 ;
        2399:  q   <=  32'b00000000000000000000000000000000 ;
        2400:  q   <=  32'b00000000000000000000000000000000 ;
        2401:  q   <=  32'b00000000000000000000000000000000 ;
        2402:  q   <=  32'b00000000000000000000000000000000 ;
        2403:  q   <=  32'b00000000000000000000000000000000 ;
        2404:  q   <=  32'b00000000000000000000000000000000 ;
        2405:  q   <=  32'b00000000000000000000000000000000 ;
        2406:  q   <=  32'b00000000000000000000000000000000 ;
        2407:  q   <=  32'b00000000000000000000000000000000 ;
        2408:  q   <=  32'b00000000000000000000000000000000 ;
        2409:  q   <=  32'b00000000000000000000000000000000 ;
        2410:  q   <=  32'b00000000000000000000000000000000 ;
        2411:  q   <=  32'b00000000000000000000000000000000 ;
        2412:  q   <=  32'b00000000000000000000000000000000 ;
        2413:  q   <=  32'b00000000000000000000000000000000 ;
        2414:  q   <=  32'b00000000000000000000000000000000 ;
        2415:  q   <=  32'b00000000000000000000000000000000 ;
        2416:  q   <=  32'b00000000000000000000000000000000 ;
        2417:  q   <=  32'b00000000000000000000000000000000 ;
        2418:  q   <=  32'b00000000000000000000000000000000 ;
        2419:  q   <=  32'b00000000000000000000000000000000 ;
        2420:  q   <=  32'b00000000000000000000000000000000 ;
        2421:  q   <=  32'b00000000000000000000000000000000 ;
        2422:  q   <=  32'b00000000000000000000000000000000 ;
        2423:  q   <=  32'b00000000000000000000000000000000 ;
        2424:  q   <=  32'b00000000000000000000000000000000 ;
        2425:  q   <=  32'b00000000000000000000000000000000 ;
        2426:  q   <=  32'b00000000000000000000000000000000 ;
        2427:  q   <=  32'b00000000000000000000000000000000 ;
        2428:  q   <=  32'b00000000000000000000000000000000 ;
        2429:  q   <=  32'b00000000000000000000000000000000 ;
        2430:  q   <=  32'b00000000000000000000000000000000 ;
        2431:  q   <=  32'b00000000000000000000000000000000 ;
        2432:  q   <=  32'b00000000000000000000000000000000 ;
        2433:  q   <=  32'b00000000000000000000000000000000 ;
        2434:  q   <=  32'b00000000000000000000000000000000 ;
        2435:  q   <=  32'b00000000000000000000000000000000 ;
        2436:  q   <=  32'b00000000000000000000000000000000 ;
        2437:  q   <=  32'b00000000000000000000000000000000 ;
        2438:  q   <=  32'b00000000000000000000000000000000 ;
        2439:  q   <=  32'b00000000000000000000000000000000 ;
        2440:  q   <=  32'b00000000000000000000000000000000 ;
        2441:  q   <=  32'b00000000000000000000000000000000 ;
        2442:  q   <=  32'b00000000000000000000000000000000 ;
        2443:  q   <=  32'b00000000000000000000000000000000 ;
        2444:  q   <=  32'b00000000000000000000000000000000 ;
        2445:  q   <=  32'b00000000000000000000000000000000 ;
        2446:  q   <=  32'b00000000000000000000000000000000 ;
        2447:  q   <=  32'b00000000000000000000000000000000 ;
        2448:  q   <=  32'b00000000000000000000000000000000 ;
        2449:  q   <=  32'b00000000000000000000000000000000 ;
        2450:  q   <=  32'b00000000000000000000000000000000 ;
        2451:  q   <=  32'b00000000000000000000000000000000 ;
        2452:  q   <=  32'b00000000000000000000000000000000 ;
        2453:  q   <=  32'b00000000000000000000000000000000 ;
        2454:  q   <=  32'b00000000000000000000000000000000 ;
        2455:  q   <=  32'b00000000000000000000000000000000 ;
        2456:  q   <=  32'b00000000000000000000000000000000 ;
        2457:  q   <=  32'b00000000000000000000000000000000 ;
        2458:  q   <=  32'b00000000000000000000000000000000 ;
        2459:  q   <=  32'b00000000000000000000000000000000 ;
        2460:  q   <=  32'b00000000000000000000000000000000 ;
        2461:  q   <=  32'b00000000000000000000000000000000 ;
        2462:  q   <=  32'b00000000000000000000000000000000 ;
        2463:  q   <=  32'b00000000000000000000000000000000 ;
        2464:  q   <=  32'b00000000000000000000000000000000 ;
        2465:  q   <=  32'b00000000000000000000000000000000 ;
        2466:  q   <=  32'b00000000000000000000000000000000 ;
        2467:  q   <=  32'b00000000000000000000000000000000 ;
        2468:  q   <=  32'b00000000000000000000000000000000 ;
        2469:  q   <=  32'b00000000000000000000000000000000 ;
        2470:  q   <=  32'b00000000000000000000000000000000 ;
        2471:  q   <=  32'b00000000000000000000000000000000 ;
        2472:  q   <=  32'b00000000000000000000000000000000 ;
        2473:  q   <=  32'b00000000000000000000000000000000 ;
        2474:  q   <=  32'b00000000000000000000000000000000 ;
        2475:  q   <=  32'b00000000000000000000000000000000 ;
        2476:  q   <=  32'b00000000000000000000000000000000 ;
        2477:  q   <=  32'b00000000000000000000000000000000 ;
        2478:  q   <=  32'b00000000000000000000000000000000 ;
        2479:  q   <=  32'b00000000000000000000000000000000 ;
        2480:  q   <=  32'b00000000000000000000000000000000 ;
        2481:  q   <=  32'b00000000000000000000000000000000 ;
        2482:  q   <=  32'b00000000000000000000000000000000 ;
        2483:  q   <=  32'b00000000000000000000000000000000 ;
        2484:  q   <=  32'b00000000000000000000000000000000 ;
        2485:  q   <=  32'b00000000000000000000000000000000 ;
        2486:  q   <=  32'b00000000000000000000000000000000 ;
        2487:  q   <=  32'b00000000000000000000000000000000 ;
        2488:  q   <=  32'b00000000000000000000000000000000 ;
        2489:  q   <=  32'b00000000000000000000000000000000 ;
        2490:  q   <=  32'b00000000000000000000000000000000 ;
        2491:  q   <=  32'b00000000000000000000000000000000 ;
        2492:  q   <=  32'b00000000000000000000000000000000 ;
        2493:  q   <=  32'b00111110011010111011100111111101 ;
        2494:  q   <=  32'b00111110111101010001101100010011 ;
        2495:  q   <=  32'b00111111001110011100010110100011 ;
        2496:  q   <=  32'b00111111011110001001011111000110 ;
        2497:  q   <=  32'b00111111100110111000001001110011 ;
        2498:  q   <=  32'b00111111101110101000011011111100 ;
        2499:  q   <=  32'b00111111110110010101100111110110 ;
        2500:  q   <=  32'b00111111111101111111101111010111 ;
        2501:  q   <=  32'b00111111111010011001001011101011 ;
        2502:  q   <=  32'b00111111110010110101000111011111 ;
        2503:  q   <=  32'b00111111101011010100000010010001 ;
        2504:  q   <=  32'b00111111100011110101111010010001 ;
        2505:  q   <=  32'b00111111011000110101011011100001 ;
        2506:  q   <=  32'b00111111001010000100110101111111 ;
        2507:  q   <=  32'b00111110110110110100000001001100 ;
        2508:  q   <=  32'b00111110010011010011011111111001 ;
        2509:  q   <=  32'b00000000000000000000000000000000 ;
        2510:  q   <=  32'b00000000000000000000000000000000 ;
        2511:  q   <=  32'b00000000000000000000000000000000 ;
        2512:  q   <=  32'b00000000000000000000000000000000 ;
        2513:  q   <=  32'b00000000000000000000000000000000 ;
        2514:  q   <=  32'b00000000000000000000000000000000 ;
        2515:  q   <=  32'b00000000000000000000000000000000 ;
        2516:  q   <=  32'b00000000000000000000000000000000 ;
        2517:  q   <=  32'b00000000000000000000000000000000 ;
        2518:  q   <=  32'b00000000000000000000000000000000 ;
        2519:  q   <=  32'b00000000000000000000000000000000 ;
        2520:  q   <=  32'b00000000000000000000000000000000 ;
        2521:  q   <=  32'b00000000000000000000000000000000 ;
        2522:  q   <=  32'b00000000000000000000000000000000 ;
        2523:  q   <=  32'b00000000000000000000000000000000 ;
        2524:  q   <=  32'b00000000000000000000000000000000 ;
        2525:  q   <=  32'b00000000000000000000000000000000 ;
        2526:  q   <=  32'b00000000000000000000000000000000 ;
        2527:  q   <=  32'b00000000000000000000000000000000 ;
        2528:  q   <=  32'b00000000000000000000000000000000 ;
        2529:  q   <=  32'b00000000000000000000000000000000 ;
        2530:  q   <=  32'b00000000000000000000000000000000 ;
        2531:  q   <=  32'b00000000000000000000000000000000 ;
        2532:  q   <=  32'b00000000000000000000000000000000 ;
        2533:  q   <=  32'b00000000000000000000000000000000 ;
        2534:  q   <=  32'b00000000000000000000000000000000 ;
        2535:  q   <=  32'b00000000000000000000000000000000 ;
        2536:  q   <=  32'b00000000000000000000000000000000 ;
        2537:  q   <=  32'b00000000000000000000000000000000 ;
        2538:  q   <=  32'b00000000000000000000000000000000 ;
        2539:  q   <=  32'b00000000000000000000000000000000 ;
        2540:  q   <=  32'b00000000000000000000000000000000 ;
        2541:  q   <=  32'b00000000000000000000000000000000 ;
        2542:  q   <=  32'b00000000000000000000000000000000 ;
        2543:  q   <=  32'b00000000000000000000000000000000 ;
        2544:  q   <=  32'b00000000000000000000000000000000 ;
        2545:  q   <=  32'b00000000000000000000000000000000 ;
        2546:  q   <=  32'b00000000000000000000000000000000 ;
        2547:  q   <=  32'b00000000000000000000000000000000 ;
        2548:  q   <=  32'b00000000000000000000000000000000 ;
        2549:  q   <=  32'b00000000000000000000000000000000 ;
        2550:  q   <=  32'b00000000000000000000000000000000 ;
        2551:  q   <=  32'b00000000000000000000000000000000 ;
        2552:  q   <=  32'b00000000000000000000000000000000 ;
        2553:  q   <=  32'b00000000000000000000000000000000 ;
        2554:  q   <=  32'b00000000000000000000000000000000 ;
        2555:  q   <=  32'b00000000000000000000000000000000 ;
        2556:  q   <=  32'b00000000000000000000000000000000 ;
        2557:  q   <=  32'b00000000000000000000000000000000 ;
        2558:  q   <=  32'b00000000000000000000000000000000 ;
        2559:  q   <=  32'b00000000000000000000000000000000 ;
        2560:  q   <=  32'b00000000000000000000000000000000 ;
        2561:  q   <=  32'b00000000000000000000000000000000 ;
        2562:  q   <=  32'b00000000000000000000000000000000 ;
        2563:  q   <=  32'b00000000000000000000000000000000 ;
        2564:  q   <=  32'b00000000000000000000000000000000 ;
        2565:  q   <=  32'b00000000000000000000000000000000 ;
        2566:  q   <=  32'b00000000000000000000000000000000 ;
        2567:  q   <=  32'b00000000000000000000000000000000 ;
        2568:  q   <=  32'b00000000000000000000000000000000 ;
        2569:  q   <=  32'b00000000000000000000000000000000 ;
        2570:  q   <=  32'b00000000000000000000000000000000 ;
        2571:  q   <=  32'b00000000000000000000000000000000 ;
        2572:  q   <=  32'b00000000000000000000000000000000 ;
        2573:  q   <=  32'b00000000000000000000000000000000 ;
        2574:  q   <=  32'b00000000000000000000000000000000 ;
        2575:  q   <=  32'b00000000000000000000000000000000 ;
        2576:  q   <=  32'b00000000000000000000000000000000 ;
        2577:  q   <=  32'b00000000000000000000000000000000 ;
        2578:  q   <=  32'b00000000000000000000000000000000 ;
        2579:  q   <=  32'b00000000000000000000000000000000 ;
        2580:  q   <=  32'b00000000000000000000000000000000 ;
        2581:  q   <=  32'b00000000000000000000000000000000 ;
        2582:  q   <=  32'b00000000000000000000000000000000 ;
        2583:  q   <=  32'b00000000000000000000000000000000 ;
        2584:  q   <=  32'b00000000000000000000000000000000 ;
        2585:  q   <=  32'b00000000000000000000000000000000 ;
        2586:  q   <=  32'b00000000000000000000000000000000 ;
        2587:  q   <=  32'b00000000000000000000000000000000 ;
        2588:  q   <=  32'b00000000000000000000000000000000 ;
        2589:  q   <=  32'b00000000000000000000000000000000 ;
        2590:  q   <=  32'b00000000000000000000000000000000 ;
        2591:  q   <=  32'b00000000000000000000000000000000 ;
        2592:  q   <=  32'b00000000000000000000000000000000 ;
        2593:  q   <=  32'b00000000000000000000000000000000 ;
        2594:  q   <=  32'b00000000000000000000000000000000 ;
        2595:  q   <=  32'b00000000000000000000000000000000 ;
        2596:  q   <=  32'b00000000000000000000000000000000 ;
        2597:  q   <=  32'b00000000000000000000000000000000 ;
        2598:  q   <=  32'b00000000000000000000000000000000 ;
        2599:  q   <=  32'b00000000000000000000000000000000 ;
        2600:  q   <=  32'b00000000000000000000000000000000 ;
        2601:  q   <=  32'b00000000000000000000000000000000 ;
        2602:  q   <=  32'b00000000000000000000000000000000 ;
        2603:  q   <=  32'b00000000000000000000000000000000 ;
        2604:  q   <=  32'b00000000000000000000000000000000 ;
        2605:  q   <=  32'b00000000000000000000000000000000 ;
        2606:  q   <=  32'b00000000000000000000000000000000 ;
        2607:  q   <=  32'b00000000000000000000000000000000 ;
        2608:  q   <=  32'b00000000000000000000000000000000 ;
        2609:  q   <=  32'b00000000000000000000000000000000 ;
        2610:  q   <=  32'b00000000000000000000000000000000 ;
        2611:  q   <=  32'b00000000000000000000000000000000 ;
        2612:  q   <=  32'b00000000000000000000000000000000 ;
        2613:  q   <=  32'b00000000000000000000000000000000 ;
        2614:  q   <=  32'b00000000000000000000000000000000 ;
        2615:  q   <=  32'b00000000000000000000000000000000 ;
        2616:  q   <=  32'b00000000000000000000000000000000 ;
        2617:  q   <=  32'b00000000000000000000000000000000 ;
        2618:  q   <=  32'b00000000000000000000000000000000 ;
        2619:  q   <=  32'b00000000000000000000000000000000 ;
        2620:  q   <=  32'b00000000000000000000000000000000 ;
        2621:  q   <=  32'b00000000000000000000000000000000 ;
        2622:  q   <=  32'b00000000000000000000000000000000 ;
        2623:  q   <=  32'b00000000000000000000000000000000 ;
        2624:  q   <=  32'b00000000000000000000000000000000 ;
        2625:  q   <=  32'b00000000000000000000000000000000 ;
        2626:  q   <=  32'b00000000000000000000000000000000 ;
        2627:  q   <=  32'b00000000000000000000000000000000 ;
        2628:  q   <=  32'b00000000000000000000000000000000 ;
        2629:  q   <=  32'b00000000000000000000000000000000 ;
        2630:  q   <=  32'b00000000000000000000000000000000 ;
        2631:  q   <=  32'b00000000000000000000000000000000 ;
        2632:  q   <=  32'b00000000000000000000000000000000 ;
        2633:  q   <=  32'b00000000000000000000000000000000 ;
        2634:  q   <=  32'b00000000000000000000000000000000 ;
        2635:  q   <=  32'b00000000000000000000000000000000 ;
        2636:  q   <=  32'b00000000000000000000000000000000 ;
        2637:  q   <=  32'b00000000000000000000000000000000 ;
        2638:  q   <=  32'b00000000000000000000000000000000 ;
        2639:  q   <=  32'b00000000000000000000000000000000 ;
        2640:  q   <=  32'b00000000000000000000000000000000 ;
        2641:  q   <=  32'b00000000000000000000000000000000 ;
        2642:  q   <=  32'b00000000000000000000000000000000 ;
        2643:  q   <=  32'b00000000000000000000000000000000 ;
        2644:  q   <=  32'b00000000000000000000000000000000 ;
        2645:  q   <=  32'b00000000000000000000000000000000 ;
        2646:  q   <=  32'b00000000000000000000000000000000 ;
        2647:  q   <=  32'b00000000000000000000000000000000 ;
        2648:  q   <=  32'b00000000000000000000000000000000 ;
        2649:  q   <=  32'b00000000000000000000000000000000 ;
        2650:  q   <=  32'b00000000000000000000000000000000 ;
        2651:  q   <=  32'b00000000000000000000000000000000 ;
        2652:  q   <=  32'b00000000000000000000000000000000 ;
        2653:  q   <=  32'b00000000000000000000000000000000 ;
        2654:  q   <=  32'b00000000000000000000000000000000 ;
        2655:  q   <=  32'b00000000000000000000000000000000 ;
        2656:  q   <=  32'b00000000000000000000000000000000 ;
        2657:  q   <=  32'b00000000000000000000000000000000 ;
        2658:  q   <=  32'b00000000000000000000000000000000 ;
        2659:  q   <=  32'b00000000000000000000000000000000 ;
        2660:  q   <=  32'b00000000000000000000000000000000 ;
        2661:  q   <=  32'b00000000000000000000000000000000 ;
        2662:  q   <=  32'b00000000000000000000000000000000 ;
        2663:  q   <=  32'b00000000000000000000000000000000 ;
        2664:  q   <=  32'b00000000000000000000000000000000 ;
        2665:  q   <=  32'b00000000000000000000000000000000 ;
        2666:  q   <=  32'b00000000000000000000000000000000 ;
        2667:  q   <=  32'b00000000000000000000000000000000 ;
        2668:  q   <=  32'b00000000000000000000000000000000 ;
        2669:  q   <=  32'b00000000000000000000000000000000 ;
        2670:  q   <=  32'b00000000000000000000000000000000 ;
        2671:  q   <=  32'b00000000000000000000000000000000 ;
        2672:  q   <=  32'b00000000000000000000000000000000 ;
        2673:  q   <=  32'b00000000000000000000000000000000 ;
        2674:  q   <=  32'b00000000000000000000000000000000 ;
        2675:  q   <=  32'b00000000000000000000000000000000 ;
        2676:  q   <=  32'b00000000000000000000000000000000 ;
        2677:  q   <=  32'b00000000000000000000000000000000 ;
        2678:  q   <=  32'b00000000000000000000000000000000 ;
        2679:  q   <=  32'b00000000000000000000000000000000 ;
        2680:  q   <=  32'b00000000000000000000000000000000 ;
        2681:  q   <=  32'b00000000000000000000000000000000 ;
        2682:  q   <=  32'b00000000000000000000000000000000 ;
        2683:  q   <=  32'b00000000000000000000000000000000 ;
        2684:  q   <=  32'b00000000000000000000000000000000 ;
        2685:  q   <=  32'b00000000000000000000000000000000 ;
        2686:  q   <=  32'b00000000000000000000000000000000 ;
        2687:  q   <=  32'b00000000000000000000000000000000 ;
        2688:  q   <=  32'b00000000000000000000000000000000 ;
        2689:  q   <=  32'b00000000000000000000000000000000 ;
        2690:  q   <=  32'b00000000000000000000000000000000 ;
        2691:  q   <=  32'b00000000000000000000000000000000 ;
        2692:  q   <=  32'b00000000000000000000000000000000 ;
        2693:  q   <=  32'b00000000000000000000000000000000 ;
        2694:  q   <=  32'b00000000000000000000000000000000 ;
        2695:  q   <=  32'b00000000000000000000000000000000 ;
        2696:  q   <=  32'b00000000000000000000000000000000 ;
        2697:  q   <=  32'b00000000000000000000000000000000 ;
        2698:  q   <=  32'b00000000000000000000000000000000 ;
        2699:  q   <=  32'b00000000000000000000000000000000 ;
        2700:  q   <=  32'b00000000000000000000000000000000 ;
        2701:  q   <=  32'b00000000000000000000000000000000 ;
        2702:  q   <=  32'b00000000000000000000000000000000 ;
        2703:  q   <=  32'b00000000000000000000000000000000 ;
        2704:  q   <=  32'b00000000000000000000000000000000 ;
        2705:  q   <=  32'b00000000000000000000000000000000 ;
        2706:  q   <=  32'b00000000000000000000000000000000 ;
        2707:  q   <=  32'b00000000000000000000000000000000 ;
        2708:  q   <=  32'b00000000000000000000000000000000 ;
        2709:  q   <=  32'b00000000000000000000000000000000 ;
        2710:  q   <=  32'b00000000000000000000000000000000 ;
        2711:  q   <=  32'b00000000000000000000000000000000 ;
        2712:  q   <=  32'b00000000000000000000000000000000 ;
        2713:  q   <=  32'b00000000000000000000000000000000 ;
        2714:  q   <=  32'b00000000000000000000000000000000 ;
        2715:  q   <=  32'b00000000000000000000000000000000 ;
        2716:  q   <=  32'b00000000000000000000000000000000 ;
        2717:  q   <=  32'b00000000000000000000000000000000 ;
        2718:  q   <=  32'b00000000000000000000000000000000 ;
        2719:  q   <=  32'b00000000000000000000000000000000 ;
        2720:  q   <=  32'b00000000000000000000000000000000 ;
        2721:  q   <=  32'b00000000000000000000000000000000 ;
        2722:  q   <=  32'b00000000000000000000000000000000 ;
        2723:  q   <=  32'b00000000000000000000000000000000 ;
        2724:  q   <=  32'b00000000000000000000000000000000 ;
        2725:  q   <=  32'b00000000000000000000000000000000 ;
        2726:  q   <=  32'b00000000000000000000000000000000 ;
        2727:  q   <=  32'b00000000000000000000000000000000 ;
        2728:  q   <=  32'b00000000000000000000000000000000 ;
        2729:  q   <=  32'b00000000000000000000000000000000 ;
        2730:  q   <=  32'b00000000000000000000000000000000 ;
        2731:  q   <=  32'b00000000000000000000000000000000 ;
        2732:  q   <=  32'b00000000000000000000000000000000 ;
        2733:  q   <=  32'b00000000000000000000000000000000 ;
        2734:  q   <=  32'b00000000000000000000000000000000 ;
        2735:  q   <=  32'b00000000000000000000000000000000 ;
        2736:  q   <=  32'b00000000000000000000000000000000 ;
        2737:  q   <=  32'b00000000000000000000000000000000 ;
        2738:  q   <=  32'b00000000000000000000000000000000 ;
        2739:  q   <=  32'b00000000000000000000000000000000 ;
        2740:  q   <=  32'b00000000000000000000000000000000 ;
        2741:  q   <=  32'b00000000000000000000000000000000 ;
        2742:  q   <=  32'b00000000000000000000000000000000 ;
        2743:  q   <=  32'b00000000000000000000000000000000 ;
        2744:  q   <=  32'b00000000000000000000000000000000 ;
        2745:  q   <=  32'b00000000000000000000000000000000 ;
        2746:  q   <=  32'b00000000000000000000000000000000 ;
        2747:  q   <=  32'b00000000000000000000000000000000 ;
        2748:  q   <=  32'b00000000000000000000000000000000 ;
        2749:  q   <=  32'b00000000000000000000000000000000 ;
        2750:  q   <=  32'b00000000000000000000000000000000 ;
        2751:  q   <=  32'b00000000000000000000000000000000 ;
        2752:  q   <=  32'b00000000000000000000000000000000 ;
        2753:  q   <=  32'b00000000000000000000000000000000 ;
        2754:  q   <=  32'b00000000000000000000000000000000 ;
        2755:  q   <=  32'b00000000000000000000000000000000 ;
        2756:  q   <=  32'b00000000000000000000000000000000 ;
        2757:  q   <=  32'b00111110001100110110100010100001 ;
        2758:  q   <=  32'b00111110110100101011100010000001 ;
        2759:  q   <=  32'b00111111001001010111111011011100 ;
        2760:  q   <=  32'b00111111011000010100001011011100 ;
        2761:  q   <=  32'b00111111100011100101010010001111 ;
        2762:  q   <=  32'b00111111101010111101100101000000 ;
        2763:  q   <=  32'b00111111110010010010111111101100 ;
        2764:  q   <=  32'b00111111111001100101100100000000 ;
        2765:  q   <=  32'b00111111111111001010101100011001 ;
        2766:  q   <=  32'b00111111110111111101101111111010 ;
        2767:  q   <=  32'b00111111110000110011100100111010 ;
        2768:  q   <=  32'b00111111101001101100001001110001 ;
        2769:  q   <=  32'b00111111100010100111011100111101 ;
        2770:  q   <=  32'b00111111010111001010111001110000 ;
        2771:  q   <=  32'b00111111001001001100010000000000 ;
        2772:  q   <=  32'b00111110110110100101110011010001 ;
        2773:  q   <=  32'b00111110010101111011001110011100 ;
        2774:  q   <=  32'b00000000000000000000000000000000 ;
        2775:  q   <=  32'b00000000000000000000000000000000 ;
        2776:  q   <=  32'b00000000000000000000000000000000 ;
        2777:  q   <=  32'b00000000000000000000000000000000 ;
        2778:  q   <=  32'b00000000000000000000000000000000 ;
        2779:  q   <=  32'b00000000000000000000000000000000 ;
        2780:  q   <=  32'b00000000000000000000000000000000 ;
        2781:  q   <=  32'b00000000000000000000000000000000 ;
        2782:  q   <=  32'b00000000000000000000000000000000 ;
        2783:  q   <=  32'b00000000000000000000000000000000 ;
        2784:  q   <=  32'b00000000000000000000000000000000 ;
        2785:  q   <=  32'b00000000000000000000000000000000 ;
        2786:  q   <=  32'b00000000000000000000000000000000 ;
        2787:  q   <=  32'b00000000000000000000000000000000 ;
        2788:  q   <=  32'b00000000000000000000000000000000 ;
        2789:  q   <=  32'b00000000000000000000000000000000 ;
        2790:  q   <=  32'b00000000000000000000000000000000 ;
        2791:  q   <=  32'b00000000000000000000000000000000 ;
        2792:  q   <=  32'b00000000000000000000000000000000 ;
        2793:  q   <=  32'b00000000000000000000000000000000 ;
        2794:  q   <=  32'b00000000000000000000000000000000 ;
        2795:  q   <=  32'b00000000000000000000000000000000 ;
        2796:  q   <=  32'b00000000000000000000000000000000 ;
        2797:  q   <=  32'b00000000000000000000000000000000 ;
        2798:  q   <=  32'b00000000000000000000000000000000 ;
        2799:  q   <=  32'b00000000000000000000000000000000 ;
        2800:  q   <=  32'b00000000000000000000000000000000 ;
        2801:  q   <=  32'b00000000000000000000000000000000 ;
        2802:  q   <=  32'b00000000000000000000000000000000 ;
        2803:  q   <=  32'b00000000000000000000000000000000 ;
        2804:  q   <=  32'b00000000000000000000000000000000 ;
        2805:  q   <=  32'b00000000000000000000000000000000 ;
        2806:  q   <=  32'b00000000000000000000000000000000 ;
        2807:  q   <=  32'b00000000000000000000000000000000 ;
        2808:  q   <=  32'b00000000000000000000000000000000 ;
        2809:  q   <=  32'b00000000000000000000000000000000 ;
        2810:  q   <=  32'b00000000000000000000000000000000 ;
        2811:  q   <=  32'b00000000000000000000000000000000 ;
        2812:  q   <=  32'b00000000000000000000000000000000 ;
        2813:  q   <=  32'b00000000000000000000000000000000 ;
        2814:  q   <=  32'b00000000000000000000000000000000 ;
        2815:  q   <=  32'b00000000000000000000000000000000 ;
        2816:  q   <=  32'b00000000000000000000000000000000 ;
        2817:  q   <=  32'b00000000000000000000000000000000 ;
        2818:  q   <=  32'b00000000000000000000000000000000 ;
        2819:  q   <=  32'b00000000000000000000000000000000 ;
        2820:  q   <=  32'b00000000000000000000000000000000 ;
        2821:  q   <=  32'b00000000000000000000000000000000 ;
        2822:  q   <=  32'b00000000000000000000000000000000 ;
        2823:  q   <=  32'b00000000000000000000000000000000 ;
        2824:  q   <=  32'b00000000000000000000000000000000 ;
        2825:  q   <=  32'b00000000000000000000000000000000 ;
        2826:  q   <=  32'b00000000000000000000000000000000 ;
        2827:  q   <=  32'b00000000000000000000000000000000 ;
        2828:  q   <=  32'b00000000000000000000000000000000 ;
        2829:  q   <=  32'b00000000000000000000000000000000 ;
        2830:  q   <=  32'b00000000000000000000000000000000 ;
        2831:  q   <=  32'b00000000000000000000000000000000 ;
        2832:  q   <=  32'b00000000000000000000000000000000 ;
        2833:  q   <=  32'b00000000000000000000000000000000 ;
        2834:  q   <=  32'b00000000000000000000000000000000 ;
        2835:  q   <=  32'b00000000000000000000000000000000 ;
        2836:  q   <=  32'b00000000000000000000000000000000 ;
        2837:  q   <=  32'b00000000000000000000000000000000 ;
        2838:  q   <=  32'b00000000000000000000000000000000 ;
        2839:  q   <=  32'b00000000000000000000000000000000 ;
        2840:  q   <=  32'b00000000000000000000000000000000 ;
        2841:  q   <=  32'b00000000000000000000000000000000 ;
        2842:  q   <=  32'b00000000000000000000000000000000 ;
        2843:  q   <=  32'b00000000000000000000000000000000 ;
        2844:  q   <=  32'b00000000000000000000000000000000 ;
        2845:  q   <=  32'b00000000000000000000000000000000 ;
        2846:  q   <=  32'b00000000000000000000000000000000 ;
        2847:  q   <=  32'b00000000000000000000000000000000 ;
        2848:  q   <=  32'b00000000000000000000000000000000 ;
        2849:  q   <=  32'b00000000000000000000000000000000 ;
        2850:  q   <=  32'b00000000000000000000000000000000 ;
        2851:  q   <=  32'b00000000000000000000000000000000 ;
        2852:  q   <=  32'b00000000000000000000000000000000 ;
        2853:  q   <=  32'b00000000000000000000000000000000 ;
        2854:  q   <=  32'b00000000000000000000000000000000 ;
        2855:  q   <=  32'b00000000000000000000000000000000 ;
        2856:  q   <=  32'b00000000000000000000000000000000 ;
        2857:  q   <=  32'b00000000000000000000000000000000 ;
        2858:  q   <=  32'b00000000000000000000000000000000 ;
        2859:  q   <=  32'b00000000000000000000000000000000 ;
        2860:  q   <=  32'b00000000000000000000000000000000 ;
        2861:  q   <=  32'b00000000000000000000000000000000 ;
        2862:  q   <=  32'b00000000000000000000000000000000 ;
        2863:  q   <=  32'b00000000000000000000000000000000 ;
        2864:  q   <=  32'b00000000000000000000000000000000 ;
        2865:  q   <=  32'b00000000000000000000000000000000 ;
        2866:  q   <=  32'b00000000000000000000000000000000 ;
        2867:  q   <=  32'b00000000000000000000000000000000 ;
        2868:  q   <=  32'b00000000000000000000000000000000 ;
        2869:  q   <=  32'b00000000000000000000000000000000 ;
        2870:  q   <=  32'b00000000000000000000000000000000 ;
        2871:  q   <=  32'b00000000000000000000000000000000 ;
        2872:  q   <=  32'b00000000000000000000000000000000 ;
        2873:  q   <=  32'b00000000000000000000000000000000 ;
        2874:  q   <=  32'b00000000000000000000000000000000 ;
        2875:  q   <=  32'b00000000000000000000000000000000 ;
        2876:  q   <=  32'b00000000000000000000000000000000 ;
        2877:  q   <=  32'b00000000000000000000000000000000 ;
        2878:  q   <=  32'b00000000000000000000000000000000 ;
        2879:  q   <=  32'b00000000000000000000000000000000 ;
        2880:  q   <=  32'b00000000000000000000000000000000 ;
        2881:  q   <=  32'b00000000000000000000000000000000 ;
        2882:  q   <=  32'b00000000000000000000000000000000 ;
        2883:  q   <=  32'b00000000000000000000000000000000 ;
        2884:  q   <=  32'b00000000000000000000000000000000 ;
        2885:  q   <=  32'b00000000000000000000000000000000 ;
        2886:  q   <=  32'b00000000000000000000000000000000 ;
        2887:  q   <=  32'b00000000000000000000000000000000 ;
        2888:  q   <=  32'b00000000000000000000000000000000 ;
        2889:  q   <=  32'b00000000000000000000000000000000 ;
        2890:  q   <=  32'b00000000000000000000000000000000 ;
        2891:  q   <=  32'b00000000000000000000000000000000 ;
        2892:  q   <=  32'b00000000000000000000000000000000 ;
        2893:  q   <=  32'b00000000000000000000000000000000 ;
        2894:  q   <=  32'b00000000000000000000000000000000 ;
        2895:  q   <=  32'b00000000000000000000000000000000 ;
        2896:  q   <=  32'b00000000000000000000000000000000 ;
        2897:  q   <=  32'b00000000000000000000000000000000 ;
        2898:  q   <=  32'b00000000000000000000000000000000 ;
        2899:  q   <=  32'b00000000000000000000000000000000 ;
        2900:  q   <=  32'b00000000000000000000000000000000 ;
        2901:  q   <=  32'b00000000000000000000000000000000 ;
        2902:  q   <=  32'b00000000000000000000000000000000 ;
        2903:  q   <=  32'b00000000000000000000000000000000 ;
        2904:  q   <=  32'b00000000000000000000000000000000 ;
        2905:  q   <=  32'b00000000000000000000000000000000 ;
        2906:  q   <=  32'b00000000000000000000000000000000 ;
        2907:  q   <=  32'b00000000000000000000000000000000 ;
        2908:  q   <=  32'b00000000000000000000000000000000 ;
        2909:  q   <=  32'b00000000000000000000000000000000 ;
        2910:  q   <=  32'b00000000000000000000000000000000 ;
        2911:  q   <=  32'b00000000000000000000000000000000 ;
        2912:  q   <=  32'b00000000000000000000000000000000 ;
        2913:  q   <=  32'b00000000000000000000000000000000 ;
        2914:  q   <=  32'b00000000000000000000000000000000 ;
        2915:  q   <=  32'b00000000000000000000000000000000 ;
        2916:  q   <=  32'b00000000000000000000000000000000 ;
        2917:  q   <=  32'b00000000000000000000000000000000 ;
        2918:  q   <=  32'b00000000000000000000000000000000 ;
        2919:  q   <=  32'b00000000000000000000000000000000 ;
        2920:  q   <=  32'b00000000000000000000000000000000 ;
        2921:  q   <=  32'b00000000000000000000000000000000 ;
        2922:  q   <=  32'b00000000000000000000000000000000 ;
        2923:  q   <=  32'b00000000000000000000000000000000 ;
        2924:  q   <=  32'b00000000000000000000000000000000 ;
        2925:  q   <=  32'b00000000000000000000000000000000 ;
        2926:  q   <=  32'b00000000000000000000000000000000 ;
        2927:  q   <=  32'b00000000000000000000000000000000 ;
        2928:  q   <=  32'b00000000000000000000000000000000 ;
        2929:  q   <=  32'b00000000000000000000000000000000 ;
        2930:  q   <=  32'b00000000000000000000000000000000 ;
        2931:  q   <=  32'b00000000000000000000000000000000 ;
        2932:  q   <=  32'b00000000000000000000000000000000 ;
        2933:  q   <=  32'b00000000000000000000000000000000 ;
        2934:  q   <=  32'b00000000000000000000000000000000 ;
        2935:  q   <=  32'b00000000000000000000000000000000 ;
        2936:  q   <=  32'b00000000000000000000000000000000 ;
        2937:  q   <=  32'b00000000000000000000000000000000 ;
        2938:  q   <=  32'b00000000000000000000000000000000 ;
        2939:  q   <=  32'b00000000000000000000000000000000 ;
        2940:  q   <=  32'b00000000000000000000000000000000 ;
        2941:  q   <=  32'b00000000000000000000000000000000 ;
        2942:  q   <=  32'b00000000000000000000000000000000 ;
        2943:  q   <=  32'b00000000000000000000000000000000 ;
        2944:  q   <=  32'b00000000000000000000000000000000 ;
        2945:  q   <=  32'b00000000000000000000000000000000 ;
        2946:  q   <=  32'b00000000000000000000000000000000 ;
        2947:  q   <=  32'b00000000000000000000000000000000 ;
        2948:  q   <=  32'b00000000000000000000000000000000 ;
        2949:  q   <=  32'b00000000000000000000000000000000 ;
        2950:  q   <=  32'b00000000000000000000000000000000 ;
        2951:  q   <=  32'b00000000000000000000000000000000 ;
        2952:  q   <=  32'b00000000000000000000000000000000 ;
        2953:  q   <=  32'b00000000000000000000000000000000 ;
        2954:  q   <=  32'b00000000000000000000000000000000 ;
        2955:  q   <=  32'b00000000000000000000000000000000 ;
        2956:  q   <=  32'b00000000000000000000000000000000 ;
        2957:  q   <=  32'b00000000000000000000000000000000 ;
        2958:  q   <=  32'b00000000000000000000000000000000 ;
        2959:  q   <=  32'b00000000000000000000000000000000 ;
        2960:  q   <=  32'b00000000000000000000000000000000 ;
        2961:  q   <=  32'b00000000000000000000000000000000 ;
        2962:  q   <=  32'b00000000000000000000000000000000 ;
        2963:  q   <=  32'b00000000000000000000000000000000 ;
        2964:  q   <=  32'b00000000000000000000000000000000 ;
        2965:  q   <=  32'b00000000000000000000000000000000 ;
        2966:  q   <=  32'b00000000000000000000000000000000 ;
        2967:  q   <=  32'b00000000000000000000000000000000 ;
        2968:  q   <=  32'b00000000000000000000000000000000 ;
        2969:  q   <=  32'b00000000000000000000000000000000 ;
        2970:  q   <=  32'b00000000000000000000000000000000 ;
        2971:  q   <=  32'b00000000000000000000000000000000 ;
        2972:  q   <=  32'b00000000000000000000000000000000 ;
        2973:  q   <=  32'b00000000000000000000000000000000 ;
        2974:  q   <=  32'b00000000000000000000000000000000 ;
        2975:  q   <=  32'b00000000000000000000000000000000 ;
        2976:  q   <=  32'b00000000000000000000000000000000 ;
        2977:  q   <=  32'b00000000000000000000000000000000 ;
        2978:  q   <=  32'b00000000000000000000000000000000 ;
        2979:  q   <=  32'b00000000000000000000000000000000 ;
        2980:  q   <=  32'b00000000000000000000000000000000 ;
        2981:  q   <=  32'b00000000000000000000000000000000 ;
        2982:  q   <=  32'b00000000000000000000000000000000 ;
        2983:  q   <=  32'b00000000000000000000000000000000 ;
        2984:  q   <=  32'b00000000000000000000000000000000 ;
        2985:  q   <=  32'b00000000000000000000000000000000 ;
        2986:  q   <=  32'b00000000000000000000000000000000 ;
        2987:  q   <=  32'b00000000000000000000000000000000 ;
        2988:  q   <=  32'b00000000000000000000000000000000 ;
        2989:  q   <=  32'b00000000000000000000000000000000 ;
        2990:  q   <=  32'b00000000000000000000000000000000 ;
        2991:  q   <=  32'b00000000000000000000000000000000 ;
        2992:  q   <=  32'b00000000000000000000000000000000 ;
        2993:  q   <=  32'b00000000000000000000000000000000 ;
        2994:  q   <=  32'b00000000000000000000000000000000 ;
        2995:  q   <=  32'b00000000000000000000000000000000 ;
        2996:  q   <=  32'b00000000000000000000000000000000 ;
        2997:  q   <=  32'b00000000000000000000000000000000 ;
        2998:  q   <=  32'b00000000000000000000000000000000 ;
        2999:  q   <=  32'b00000000000000000000000000000000 ;
        3000:  q   <=  32'b00000000000000000000000000000000 ;
        3001:  q   <=  32'b00000000000000000000000000000000 ;
        3002:  q   <=  32'b00000000000000000000000000000000 ;
        3003:  q   <=  32'b00000000000000000000000000000000 ;
        3004:  q   <=  32'b00000000000000000000000000000000 ;
        3005:  q   <=  32'b00000000000000000000000000000000 ;
        3006:  q   <=  32'b00000000000000000000000000000000 ;
        3007:  q   <=  32'b00000000000000000000000000000000 ;
        3008:  q   <=  32'b00000000000000000000000000000000 ;
        3009:  q   <=  32'b00000000000000000000000000000000 ;
        3010:  q   <=  32'b00000000000000000000000000000000 ;
        3011:  q   <=  32'b00000000000000000000000000000000 ;
        3012:  q   <=  32'b00000000000000000000000000000000 ;
        3013:  q   <=  32'b00000000000000000000000000000000 ;
        3014:  q   <=  32'b00000000000000000000000000000000 ;
        3015:  q   <=  32'b00000000000000000000000000000000 ;
        3016:  q   <=  32'b00000000000000000000000000000000 ;
        3017:  q   <=  32'b00000000000000000000000000000000 ;
        3018:  q   <=  32'b00000000000000000000000000000000 ;
        3019:  q   <=  32'b00000000000000000000000000000000 ;
        3020:  q   <=  32'b00000000000000000000000000000000 ;
        3021:  q   <=  32'b00111100110101010011100110001000 ;
        3022:  q   <=  32'b00111110100000001001000000010101 ;
        3023:  q   <=  32'b00111110111100110001101100010111 ;
        3024:  q   <=  32'b00111111001100100111101100011100 ;
        3025:  q   <=  32'b00111111011010110001000110000101 ;
        3026:  q   <=  32'b00111111100100011010100011000111 ;
        3027:  q   <=  32'b00111111101011011001110111111111 ;
        3028:  q   <=  32'b00111111110010010110100011001011 ;
        3029:  q   <=  32'b00111111111001010000100110001100 ;
        3030:  q   <=  32'b00111111111111110111111101011111 ;
        3031:  q   <=  32'b00111111111001000011000110011001 ;
        3032:  q   <=  32'b00111111110010010000110011000100 ;
        3033:  q   <=  32'b00111111101011100001000010000101 ;
        3034:  q   <=  32'b00111111100100110011110010000000 ;
        3035:  q   <=  32'b00111111011100010010000010111010 ;
        3036:  q   <=  32'b00111111001111000001011110000101 ;
        3037:  q   <=  32'b00111111000001110101110010110001 ;
        3038:  q   <=  32'b00111110101001011101111100100010 ;
        3039:  q   <=  32'b00111101111101100111101111010110 ;
        3040:  q   <=  32'b00000000000000000000000000000000 ;
        3041:  q   <=  32'b00000000000000000000000000000000 ;
        3042:  q   <=  32'b00000000000000000000000000000000 ;
        3043:  q   <=  32'b00000000000000000000000000000000 ;
        3044:  q   <=  32'b00000000000000000000000000000000 ;
        3045:  q   <=  32'b00000000000000000000000000000000 ;
        3046:  q   <=  32'b00000000000000000000000000000000 ;
        3047:  q   <=  32'b00000000000000000000000000000000 ;
        3048:  q   <=  32'b00000000000000000000000000000000 ;
        3049:  q   <=  32'b00000000000000000000000000000000 ;
        3050:  q   <=  32'b00000000000000000000000000000000 ;
        3051:  q   <=  32'b00000000000000000000000000000000 ;
        3052:  q   <=  32'b00000000000000000000000000000000 ;
        3053:  q   <=  32'b00000000000000000000000000000000 ;
        3054:  q   <=  32'b00000000000000000000000000000000 ;
        3055:  q   <=  32'b00000000000000000000000000000000 ;
        3056:  q   <=  32'b00000000000000000000000000000000 ;
        3057:  q   <=  32'b00000000000000000000000000000000 ;
        3058:  q   <=  32'b00000000000000000000000000000000 ;
        3059:  q   <=  32'b00000000000000000000000000000000 ;
        3060:  q   <=  32'b00000000000000000000000000000000 ;
        3061:  q   <=  32'b00000000000000000000000000000000 ;
        3062:  q   <=  32'b00000000000000000000000000000000 ;
        3063:  q   <=  32'b00000000000000000000000000000000 ;
        3064:  q   <=  32'b00000000000000000000000000000000 ;
        3065:  q   <=  32'b00000000000000000000000000000000 ;
        3066:  q   <=  32'b00000000000000000000000000000000 ;
        3067:  q   <=  32'b00000000000000000000000000000000 ;
        3068:  q   <=  32'b00000000000000000000000000000000 ;
        3069:  q   <=  32'b00000000000000000000000000000000 ;
        3070:  q   <=  32'b00000000000000000000000000000000 ;
        3071:  q   <=  32'b00000000000000000000000000000000 ;
        3072:  q   <=  32'b00000000000000000000000000000000 ;
        3073:  q   <=  32'b00000000000000000000000000000000 ;
        3074:  q   <=  32'b00000000000000000000000000000000 ;
        3075:  q   <=  32'b00000000000000000000000000000000 ;
        3076:  q   <=  32'b00000000000000000000000000000000 ;
        3077:  q   <=  32'b00000000000000000000000000000000 ;
        3078:  q   <=  32'b00000000000000000000000000000000 ;
        3079:  q   <=  32'b00000000000000000000000000000000 ;
        3080:  q   <=  32'b00000000000000000000000000000000 ;
        3081:  q   <=  32'b00000000000000000000000000000000 ;
        3082:  q   <=  32'b00000000000000000000000000000000 ;
        3083:  q   <=  32'b00000000000000000000000000000000 ;
        3084:  q   <=  32'b00000000000000000000000000000000 ;
        3085:  q   <=  32'b00000000000000000000000000000000 ;
        3086:  q   <=  32'b00000000000000000000000000000000 ;
        3087:  q   <=  32'b00000000000000000000000000000000 ;
        3088:  q   <=  32'b00000000000000000000000000000000 ;
        3089:  q   <=  32'b00000000000000000000000000000000 ;
        3090:  q   <=  32'b00000000000000000000000000000000 ;
        3091:  q   <=  32'b00000000000000000000000000000000 ;
        3092:  q   <=  32'b00000000000000000000000000000000 ;
        3093:  q   <=  32'b00000000000000000000000000000000 ;
        3094:  q   <=  32'b00000000000000000000000000000000 ;
        3095:  q   <=  32'b00000000000000000000000000000000 ;
        3096:  q   <=  32'b00000000000000000000000000000000 ;
        3097:  q   <=  32'b00000000000000000000000000000000 ;
        3098:  q   <=  32'b00000000000000000000000000000000 ;
        3099:  q   <=  32'b00000000000000000000000000000000 ;
        3100:  q   <=  32'b00000000000000000000000000000000 ;
        3101:  q   <=  32'b00000000000000000000000000000000 ;
        3102:  q   <=  32'b00000000000000000000000000000000 ;
        3103:  q   <=  32'b00000000000000000000000000000000 ;
        3104:  q   <=  32'b00000000000000000000000000000000 ;
        3105:  q   <=  32'b00000000000000000000000000000000 ;
        3106:  q   <=  32'b00000000000000000000000000000000 ;
        3107:  q   <=  32'b00000000000000000000000000000000 ;
        3108:  q   <=  32'b00000000000000000000000000000000 ;
        3109:  q   <=  32'b00000000000000000000000000000000 ;
        3110:  q   <=  32'b00000000000000000000000000000000 ;
        3111:  q   <=  32'b00000000000000000000000000000000 ;
        3112:  q   <=  32'b00000000000000000000000000000000 ;
        3113:  q   <=  32'b00000000000000000000000000000000 ;
        3114:  q   <=  32'b00000000000000000000000000000000 ;
        3115:  q   <=  32'b00000000000000000000000000000000 ;
        3116:  q   <=  32'b00000000000000000000000000000000 ;
        3117:  q   <=  32'b00000000000000000000000000000000 ;
        3118:  q   <=  32'b00000000000000000000000000000000 ;
        3119:  q   <=  32'b00000000000000000000000000000000 ;
        3120:  q   <=  32'b00000000000000000000000000000000 ;
        3121:  q   <=  32'b00000000000000000000000000000000 ;
        3122:  q   <=  32'b00000000000000000000000000000000 ;
        3123:  q   <=  32'b00000000000000000000000000000000 ;
        3124:  q   <=  32'b00000000000000000000000000000000 ;
        3125:  q   <=  32'b00000000000000000000000000000000 ;
        3126:  q   <=  32'b00000000000000000000000000000000 ;
        3127:  q   <=  32'b00000000000000000000000000000000 ;
        3128:  q   <=  32'b00000000000000000000000000000000 ;
        3129:  q   <=  32'b00000000000000000000000000000000 ;
        3130:  q   <=  32'b00000000000000000000000000000000 ;
        3131:  q   <=  32'b00000000000000000000000000000000 ;
        3132:  q   <=  32'b00000000000000000000000000000000 ;
        3133:  q   <=  32'b00000000000000000000000000000000 ;
        3134:  q   <=  32'b00000000000000000000000000000000 ;
        3135:  q   <=  32'b00000000000000000000000000000000 ;
        3136:  q   <=  32'b00000000000000000000000000000000 ;
        3137:  q   <=  32'b00000000000000000000000000000000 ;
        3138:  q   <=  32'b00000000000000000000000000000000 ;
        3139:  q   <=  32'b00000000000000000000000000000000 ;
        3140:  q   <=  32'b00000000000000000000000000000000 ;
        3141:  q   <=  32'b00000000000000000000000000000000 ;
        3142:  q   <=  32'b00000000000000000000000000000000 ;
        3143:  q   <=  32'b00000000000000000000000000000000 ;
        3144:  q   <=  32'b00000000000000000000000000000000 ;
        3145:  q   <=  32'b00000000000000000000000000000000 ;
        3146:  q   <=  32'b00000000000000000000000000000000 ;
        3147:  q   <=  32'b00000000000000000000000000000000 ;
        3148:  q   <=  32'b00000000000000000000000000000000 ;
        3149:  q   <=  32'b00000000000000000000000000000000 ;
        3150:  q   <=  32'b00000000000000000000000000000000 ;
        3151:  q   <=  32'b00000000000000000000000000000000 ;
        3152:  q   <=  32'b00000000000000000000000000000000 ;
        3153:  q   <=  32'b00000000000000000000000000000000 ;
        3154:  q   <=  32'b00000000000000000000000000000000 ;
        3155:  q   <=  32'b00000000000000000000000000000000 ;
        3156:  q   <=  32'b00000000000000000000000000000000 ;
        3157:  q   <=  32'b00000000000000000000000000000000 ;
        3158:  q   <=  32'b00000000000000000000000000000000 ;
        3159:  q   <=  32'b00000000000000000000000000000000 ;
        3160:  q   <=  32'b00000000000000000000000000000000 ;
        3161:  q   <=  32'b00000000000000000000000000000000 ;
        3162:  q   <=  32'b00000000000000000000000000000000 ;
        3163:  q   <=  32'b00000000000000000000000000000000 ;
        3164:  q   <=  32'b00000000000000000000000000000000 ;
        3165:  q   <=  32'b00000000000000000000000000000000 ;
        3166:  q   <=  32'b00000000000000000000000000000000 ;
        3167:  q   <=  32'b00000000000000000000000000000000 ;
        3168:  q   <=  32'b00000000000000000000000000000000 ;
        3169:  q   <=  32'b00000000000000000000000000000000 ;
        3170:  q   <=  32'b00000000000000000000000000000000 ;
        3171:  q   <=  32'b00000000000000000000000000000000 ;
        3172:  q   <=  32'b00000000000000000000000000000000 ;
        3173:  q   <=  32'b00000000000000000000000000000000 ;
        3174:  q   <=  32'b00000000000000000000000000000000 ;
        3175:  q   <=  32'b00000000000000000000000000000000 ;
        3176:  q   <=  32'b00000000000000000000000000000000 ;
        3177:  q   <=  32'b00000000000000000000000000000000 ;
        3178:  q   <=  32'b00000000000000000000000000000000 ;
        3179:  q   <=  32'b00000000000000000000000000000000 ;
        3180:  q   <=  32'b00000000000000000000000000000000 ;
        3181:  q   <=  32'b00000000000000000000000000000000 ;
        3182:  q   <=  32'b00000000000000000000000000000000 ;
        3183:  q   <=  32'b00000000000000000000000000000000 ;
        3184:  q   <=  32'b00000000000000000000000000000000 ;
        3185:  q   <=  32'b00000000000000000000000000000000 ;
        3186:  q   <=  32'b00000000000000000000000000000000 ;
        3187:  q   <=  32'b00000000000000000000000000000000 ;
        3188:  q   <=  32'b00000000000000000000000000000000 ;
        3189:  q   <=  32'b00000000000000000000000000000000 ;
        3190:  q   <=  32'b00000000000000000000000000000000 ;
        3191:  q   <=  32'b00000000000000000000000000000000 ;
        3192:  q   <=  32'b00000000000000000000000000000000 ;
        3193:  q   <=  32'b00000000000000000000000000000000 ;
        3194:  q   <=  32'b00000000000000000000000000000000 ;
        3195:  q   <=  32'b00000000000000000000000000000000 ;
        3196:  q   <=  32'b00000000000000000000000000000000 ;
        3197:  q   <=  32'b00000000000000000000000000000000 ;
        3198:  q   <=  32'b00000000000000000000000000000000 ;
        3199:  q   <=  32'b00000000000000000000000000000000 ;
        3200:  q   <=  32'b00000000000000000000000000000000 ;
        3201:  q   <=  32'b00000000000000000000000000000000 ;
        3202:  q   <=  32'b00000000000000000000000000000000 ;
        3203:  q   <=  32'b00000000000000000000000000000000 ;
        3204:  q   <=  32'b00000000000000000000000000000000 ;
        3205:  q   <=  32'b00000000000000000000000000000000 ;
        3206:  q   <=  32'b00000000000000000000000000000000 ;
        3207:  q   <=  32'b00000000000000000000000000000000 ;
        3208:  q   <=  32'b00000000000000000000000000000000 ;
        3209:  q   <=  32'b00000000000000000000000000000000 ;
        3210:  q   <=  32'b00000000000000000000000000000000 ;
        3211:  q   <=  32'b00000000000000000000000000000000 ;
        3212:  q   <=  32'b00000000000000000000000000000000 ;
        3213:  q   <=  32'b00000000000000000000000000000000 ;
        3214:  q   <=  32'b00000000000000000000000000000000 ;
        3215:  q   <=  32'b00000000000000000000000000000000 ;
        3216:  q   <=  32'b00000000000000000000000000000000 ;
        3217:  q   <=  32'b00000000000000000000000000000000 ;
        3218:  q   <=  32'b00000000000000000000000000000000 ;
        3219:  q   <=  32'b00000000000000000000000000000000 ;
        3220:  q   <=  32'b00000000000000000000000000000000 ;
        3221:  q   <=  32'b00000000000000000000000000000000 ;
        3222:  q   <=  32'b00000000000000000000000000000000 ;
        3223:  q   <=  32'b00000000000000000000000000000000 ;
        3224:  q   <=  32'b00000000000000000000000000000000 ;
        3225:  q   <=  32'b00000000000000000000000000000000 ;
        3226:  q   <=  32'b00000000000000000000000000000000 ;
        3227:  q   <=  32'b00000000000000000000000000000000 ;
        3228:  q   <=  32'b00000000000000000000000000000000 ;
        3229:  q   <=  32'b00000000000000000000000000000000 ;
        3230:  q   <=  32'b00000000000000000000000000000000 ;
        3231:  q   <=  32'b00000000000000000000000000000000 ;
        3232:  q   <=  32'b00000000000000000000000000000000 ;
        3233:  q   <=  32'b00000000000000000000000000000000 ;
        3234:  q   <=  32'b00000000000000000000000000000000 ;
        3235:  q   <=  32'b00000000000000000000000000000000 ;
        3236:  q   <=  32'b00000000000000000000000000000000 ;
        3237:  q   <=  32'b00000000000000000000000000000000 ;
        3238:  q   <=  32'b00000000000000000000000000000000 ;
        3239:  q   <=  32'b00000000000000000000000000000000 ;
        3240:  q   <=  32'b00000000000000000000000000000000 ;
        3241:  q   <=  32'b00000000000000000000000000000000 ;
        3242:  q   <=  32'b00000000000000000000000000000000 ;
        3243:  q   <=  32'b00000000000000000000000000000000 ;
        3244:  q   <=  32'b00000000000000000000000000000000 ;
        3245:  q   <=  32'b00000000000000000000000000000000 ;
        3246:  q   <=  32'b00000000000000000000000000000000 ;
        3247:  q   <=  32'b00000000000000000000000000000000 ;
        3248:  q   <=  32'b00000000000000000000000000000000 ;
        3249:  q   <=  32'b00000000000000000000000000000000 ;
        3250:  q   <=  32'b00000000000000000000000000000000 ;
        3251:  q   <=  32'b00000000000000000000000000000000 ;
        3252:  q   <=  32'b00000000000000000000000000000000 ;
        3253:  q   <=  32'b00000000000000000000000000000000 ;
        3254:  q   <=  32'b00000000000000000000000000000000 ;
        3255:  q   <=  32'b00000000000000000000000000000000 ;
        3256:  q   <=  32'b00000000000000000000000000000000 ;
        3257:  q   <=  32'b00000000000000000000000000000000 ;
        3258:  q   <=  32'b00000000000000000000000000000000 ;
        3259:  q   <=  32'b00000000000000000000000000000000 ;
        3260:  q   <=  32'b00000000000000000000000000000000 ;
        3261:  q   <=  32'b00000000000000000000000000000000 ;
        3262:  q   <=  32'b00000000000000000000000000000000 ;
        3263:  q   <=  32'b00000000000000000000000000000000 ;
        3264:  q   <=  32'b00000000000000000000000000000000 ;
        3265:  q   <=  32'b00000000000000000000000000000000 ;
        3266:  q   <=  32'b00000000000000000000000000000000 ;
        3267:  q   <=  32'b00000000000000000000000000000000 ;
        3268:  q   <=  32'b00000000000000000000000000000000 ;
        3269:  q   <=  32'b00000000000000000000000000000000 ;
        3270:  q   <=  32'b00000000000000000000000000000000 ;
        3271:  q   <=  32'b00000000000000000000000000000000 ;
        3272:  q   <=  32'b00000000000000000000000000000000 ;
        3273:  q   <=  32'b00000000000000000000000000000000 ;
        3274:  q   <=  32'b00000000000000000000000000000000 ;
        3275:  q   <=  32'b00000000000000000000000000000000 ;
        3276:  q   <=  32'b00000000000000000000000000000000 ;
        3277:  q   <=  32'b00000000000000000000000000000000 ;
        3278:  q   <=  32'b00000000000000000000000000000000 ;
        3279:  q   <=  32'b00000000000000000000000000000000 ;
        3280:  q   <=  32'b00000000000000000000000000000000 ;
        3281:  q   <=  32'b00000000000000000000000000000000 ;
        3282:  q   <=  32'b00000000000000000000000000000000 ;
        3283:  q   <=  32'b00000000000000000000000000000000 ;
        3284:  q   <=  32'b00000000000000000000000000000000 ;
        3285:  q   <=  32'b00000000000000000000000000000000 ;
        3286:  q   <=  32'b00111011100000001010000011011011 ;
        3287:  q   <=  32'b00111110010111100111001100110111 ;
        3288:  q   <=  32'b00111110110110111100110011101110 ;
        3289:  q   <=  32'b00111111001000111101111011110101 ;
        3290:  q   <=  32'b00111111010110011000011011111110 ;
        3291:  q   <=  32'b00111111100001110110111110100010 ;
        3292:  q   <=  32'b00111111101000011111010000111101 ;
        3293:  q   <=  32'b00111111101111000101000110100111 ;
        3294:  q   <=  32'b00111111110101101000100000110111 ;
        3295:  q   <=  32'b00111111111100001001100001000010 ;
        3296:  q   <=  32'b00111111111101010111110111100001 ;
        3297:  q   <=  32'b00111111110110111011100111100010 ;
        3298:  q   <=  32'b00111111110000100001101101101101 ;
        3299:  q   <=  32'b00111111101010001010001000101110 ;
        3300:  q   <=  32'b00111111100011110100110111010111 ;
        3301:  q   <=  32'b00111111011011000011110000101110 ;
        3302:  q   <=  32'b00111111001110100010010100111101 ;
        3303:  q   <=  32'b00111111000010000101011000111111 ;
        3304:  q   <=  32'b00111110101011011001110100110011 ;
        3305:  q   <=  32'b00111110000101100011011011001111 ;
        3306:  q   <=  32'b00000000000000000000000000000000 ;
        3307:  q   <=  32'b00000000000000000000000000000000 ;
        3308:  q   <=  32'b00000000000000000000000000000000 ;
        3309:  q   <=  32'b00000000000000000000000000000000 ;
        3310:  q   <=  32'b00000000000000000000000000000000 ;
        3311:  q   <=  32'b00000000000000000000000000000000 ;
        3312:  q   <=  32'b00000000000000000000000000000000 ;
        3313:  q   <=  32'b00000000000000000000000000000000 ;
        3314:  q   <=  32'b00000000000000000000000000000000 ;
        3315:  q   <=  32'b00000000000000000000000000000000 ;
        3316:  q   <=  32'b00000000000000000000000000000000 ;
        3317:  q   <=  32'b00000000000000000000000000000000 ;
        3318:  q   <=  32'b00000000000000000000000000000000 ;
        3319:  q   <=  32'b00000000000000000000000000000000 ;
        3320:  q   <=  32'b00000000000000000000000000000000 ;
        3321:  q   <=  32'b00000000000000000000000000000000 ;
        3322:  q   <=  32'b00000000000000000000000000000000 ;
        3323:  q   <=  32'b00000000000000000000000000000000 ;
        3324:  q   <=  32'b00000000000000000000000000000000 ;
        3325:  q   <=  32'b00000000000000000000000000000000 ;
        3326:  q   <=  32'b00000000000000000000000000000000 ;
        3327:  q   <=  32'b00000000000000000000000000000000 ;
        3328:  q   <=  32'b00000000000000000000000000000000 ;
        3329:  q   <=  32'b00000000000000000000000000000000 ;
        3330:  q   <=  32'b00000000000000000000000000000000 ;
        3331:  q   <=  32'b00000000000000000000000000000000 ;
        3332:  q   <=  32'b00000000000000000000000000000000 ;
        3333:  q   <=  32'b00000000000000000000000000000000 ;
        3334:  q   <=  32'b00000000000000000000000000000000 ;
        3335:  q   <=  32'b00000000000000000000000000000000 ;
        3336:  q   <=  32'b00000000000000000000000000000000 ;
        3337:  q   <=  32'b00000000000000000000000000000000 ;
        3338:  q   <=  32'b00000000000000000000000000000000 ;
        3339:  q   <=  32'b00000000000000000000000000000000 ;
        3340:  q   <=  32'b00000000000000000000000000000000 ;
        3341:  q   <=  32'b00000000000000000000000000000000 ;
        3342:  q   <=  32'b00000000000000000000000000000000 ;
        3343:  q   <=  32'b00000000000000000000000000000000 ;
        3344:  q   <=  32'b00000000000000000000000000000000 ;
        3345:  q   <=  32'b00000000000000000000000000000000 ;
        3346:  q   <=  32'b00000000000000000000000000000000 ;
        3347:  q   <=  32'b00000000000000000000000000000000 ;
        3348:  q   <=  32'b00000000000000000000000000000000 ;
        3349:  q   <=  32'b00000000000000000000000000000000 ;
        3350:  q   <=  32'b00000000000000000000000000000000 ;
        3351:  q   <=  32'b00000000000000000000000000000000 ;
        3352:  q   <=  32'b00000000000000000000000000000000 ;
        3353:  q   <=  32'b00000000000000000000000000000000 ;
        3354:  q   <=  32'b00000000000000000000000000000000 ;
        3355:  q   <=  32'b00000000000000000000000000000000 ;
        3356:  q   <=  32'b00000000000000000000000000000000 ;
        3357:  q   <=  32'b00000000000000000000000000000000 ;
        3358:  q   <=  32'b00000000000000000000000000000000 ;
        3359:  q   <=  32'b00000000000000000000000000000000 ;
        3360:  q   <=  32'b00000000000000000000000000000000 ;
        3361:  q   <=  32'b00000000000000000000000000000000 ;
        3362:  q   <=  32'b00000000000000000000000000000000 ;
        3363:  q   <=  32'b00000000000000000000000000000000 ;
        3364:  q   <=  32'b00000000000000000000000000000000 ;
        3365:  q   <=  32'b00000000000000000000000000000000 ;
        3366:  q   <=  32'b00000000000000000000000000000000 ;
        3367:  q   <=  32'b00000000000000000000000000000000 ;
        3368:  q   <=  32'b00000000000000000000000000000000 ;
        3369:  q   <=  32'b00000000000000000000000000000000 ;
        3370:  q   <=  32'b00000000000000000000000000000000 ;
        3371:  q   <=  32'b00000000000000000000000000000000 ;
        3372:  q   <=  32'b00000000000000000000000000000000 ;
        3373:  q   <=  32'b00000000000000000000000000000000 ;
        3374:  q   <=  32'b00000000000000000000000000000000 ;
        3375:  q   <=  32'b00000000000000000000000000000000 ;
        3376:  q   <=  32'b00000000000000000000000000000000 ;
        3377:  q   <=  32'b00000000000000000000000000000000 ;
        3378:  q   <=  32'b00000000000000000000000000000000 ;
        3379:  q   <=  32'b00000000000000000000000000000000 ;
        3380:  q   <=  32'b00000000000000000000000000000000 ;
        3381:  q   <=  32'b00000000000000000000000000000000 ;
        3382:  q   <=  32'b00000000000000000000000000000000 ;
        3383:  q   <=  32'b00000000000000000000000000000000 ;
        3384:  q   <=  32'b00000000000000000000000000000000 ;
        3385:  q   <=  32'b00000000000000000000000000000000 ;
        3386:  q   <=  32'b00000000000000000000000000000000 ;
        3387:  q   <=  32'b00000000000000000000000000000000 ;
        3388:  q   <=  32'b00000000000000000000000000000000 ;
        3389:  q   <=  32'b00000000000000000000000000000000 ;
        3390:  q   <=  32'b00000000000000000000000000000000 ;
        3391:  q   <=  32'b00000000000000000000000000000000 ;
        3392:  q   <=  32'b00000000000000000000000000000000 ;
        3393:  q   <=  32'b00000000000000000000000000000000 ;
        3394:  q   <=  32'b00000000000000000000000000000000 ;
        3395:  q   <=  32'b00000000000000000000000000000000 ;
        3396:  q   <=  32'b00000000000000000000000000000000 ;
        3397:  q   <=  32'b00000000000000000000000000000000 ;
        3398:  q   <=  32'b00000000000000000000000000000000 ;
        3399:  q   <=  32'b00000000000000000000000000000000 ;
        3400:  q   <=  32'b00000000000000000000000000000000 ;
        3401:  q   <=  32'b00000000000000000000000000000000 ;
        3402:  q   <=  32'b00000000000000000000000000000000 ;
        3403:  q   <=  32'b00000000000000000000000000000000 ;
        3404:  q   <=  32'b00000000000000000000000000000000 ;
        3405:  q   <=  32'b00000000000000000000000000000000 ;
        3406:  q   <=  32'b00000000000000000000000000000000 ;
        3407:  q   <=  32'b00000000000000000000000000000000 ;
        3408:  q   <=  32'b00000000000000000000000000000000 ;
        3409:  q   <=  32'b00000000000000000000000000000000 ;
        3410:  q   <=  32'b00000000000000000000000000000000 ;
        3411:  q   <=  32'b00000000000000000000000000000000 ;
        3412:  q   <=  32'b00000000000000000000000000000000 ;
        3413:  q   <=  32'b00000000000000000000000000000000 ;
        3414:  q   <=  32'b00000000000000000000000000000000 ;
        3415:  q   <=  32'b00000000000000000000000000000000 ;
        3416:  q   <=  32'b00000000000000000000000000000000 ;
        3417:  q   <=  32'b00000000000000000000000000000000 ;
        3418:  q   <=  32'b00000000000000000000000000000000 ;
        3419:  q   <=  32'b00000000000000000000000000000000 ;
        3420:  q   <=  32'b00000000000000000000000000000000 ;
        3421:  q   <=  32'b00000000000000000000000000000000 ;
        3422:  q   <=  32'b00000000000000000000000000000000 ;
        3423:  q   <=  32'b00000000000000000000000000000000 ;
        3424:  q   <=  32'b00000000000000000000000000000000 ;
        3425:  q   <=  32'b00000000000000000000000000000000 ;
        3426:  q   <=  32'b00000000000000000000000000000000 ;
        3427:  q   <=  32'b00000000000000000000000000000000 ;
        3428:  q   <=  32'b00000000000000000000000000000000 ;
        3429:  q   <=  32'b00000000000000000000000000000000 ;
        3430:  q   <=  32'b00000000000000000000000000000000 ;
        3431:  q   <=  32'b00000000000000000000000000000000 ;
        3432:  q   <=  32'b00000000000000000000000000000000 ;
        3433:  q   <=  32'b00000000000000000000000000000000 ;
        3434:  q   <=  32'b00000000000000000000000000000000 ;
        3435:  q   <=  32'b00000000000000000000000000000000 ;
        3436:  q   <=  32'b00000000000000000000000000000000 ;
        3437:  q   <=  32'b00000000000000000000000000000000 ;
        3438:  q   <=  32'b00000000000000000000000000000000 ;
        3439:  q   <=  32'b00000000000000000000000000000000 ;
        3440:  q   <=  32'b00000000000000000000000000000000 ;
        3441:  q   <=  32'b00000000000000000000000000000000 ;
        3442:  q   <=  32'b00000000000000000000000000000000 ;
        3443:  q   <=  32'b00000000000000000000000000000000 ;
        3444:  q   <=  32'b00000000000000000000000000000000 ;
        3445:  q   <=  32'b00000000000000000000000000000000 ;
        3446:  q   <=  32'b00000000000000000000000000000000 ;
        3447:  q   <=  32'b00000000000000000000000000000000 ;
        3448:  q   <=  32'b00000000000000000000000000000000 ;
        3449:  q   <=  32'b00000000000000000000000000000000 ;
        3450:  q   <=  32'b00000000000000000000000000000000 ;
        3451:  q   <=  32'b00000000000000000000000000000000 ;
        3452:  q   <=  32'b00000000000000000000000000000000 ;
        3453:  q   <=  32'b00000000000000000000000000000000 ;
        3454:  q   <=  32'b00000000000000000000000000000000 ;
        3455:  q   <=  32'b00000000000000000000000000000000 ;
        3456:  q   <=  32'b00000000000000000000000000000000 ;
        3457:  q   <=  32'b00000000000000000000000000000000 ;
        3458:  q   <=  32'b00000000000000000000000000000000 ;
        3459:  q   <=  32'b00000000000000000000000000000000 ;
        3460:  q   <=  32'b00000000000000000000000000000000 ;
        3461:  q   <=  32'b00000000000000000000000000000000 ;
        3462:  q   <=  32'b00000000000000000000000000000000 ;
        3463:  q   <=  32'b00000000000000000000000000000000 ;
        3464:  q   <=  32'b00000000000000000000000000000000 ;
        3465:  q   <=  32'b00000000000000000000000000000000 ;
        3466:  q   <=  32'b00000000000000000000000000000000 ;
        3467:  q   <=  32'b00000000000000000000000000000000 ;
        3468:  q   <=  32'b00000000000000000000000000000000 ;
        3469:  q   <=  32'b00000000000000000000000000000000 ;
        3470:  q   <=  32'b00000000000000000000000000000000 ;
        3471:  q   <=  32'b00000000000000000000000000000000 ;
        3472:  q   <=  32'b00000000000000000000000000000000 ;
        3473:  q   <=  32'b00000000000000000000000000000000 ;
        3474:  q   <=  32'b00000000000000000000000000000000 ;
        3475:  q   <=  32'b00000000000000000000000000000000 ;
        3476:  q   <=  32'b00000000000000000000000000000000 ;
        3477:  q   <=  32'b00000000000000000000000000000000 ;
        3478:  q   <=  32'b00000000000000000000000000000000 ;
        3479:  q   <=  32'b00000000000000000000000000000000 ;
        3480:  q   <=  32'b00000000000000000000000000000000 ;
        3481:  q   <=  32'b00000000000000000000000000000000 ;
        3482:  q   <=  32'b00000000000000000000000000000000 ;
        3483:  q   <=  32'b00000000000000000000000000000000 ;
        3484:  q   <=  32'b00000000000000000000000000000000 ;
        3485:  q   <=  32'b00000000000000000000000000000000 ;
        3486:  q   <=  32'b00000000000000000000000000000000 ;
        3487:  q   <=  32'b00000000000000000000000000000000 ;
        3488:  q   <=  32'b00000000000000000000000000000000 ;
        3489:  q   <=  32'b00000000000000000000000000000000 ;
        3490:  q   <=  32'b00000000000000000000000000000000 ;
        3491:  q   <=  32'b00000000000000000000000000000000 ;
        3492:  q   <=  32'b00000000000000000000000000000000 ;
        3493:  q   <=  32'b00000000000000000000000000000000 ;
        3494:  q   <=  32'b00000000000000000000000000000000 ;
        3495:  q   <=  32'b00000000000000000000000000000000 ;
        3496:  q   <=  32'b00000000000000000000000000000000 ;
        3497:  q   <=  32'b00000000000000000000000000000000 ;
        3498:  q   <=  32'b00000000000000000000000000000000 ;
        3499:  q   <=  32'b00000000000000000000000000000000 ;
        3500:  q   <=  32'b00000000000000000000000000000000 ;
        3501:  q   <=  32'b00000000000000000000000000000000 ;
        3502:  q   <=  32'b00000000000000000000000000000000 ;
        3503:  q   <=  32'b00000000000000000000000000000000 ;
        3504:  q   <=  32'b00000000000000000000000000000000 ;
        3505:  q   <=  32'b00000000000000000000000000000000 ;
        3506:  q   <=  32'b00000000000000000000000000000000 ;
        3507:  q   <=  32'b00000000000000000000000000000000 ;
        3508:  q   <=  32'b00000000000000000000000000000000 ;
        3509:  q   <=  32'b00000000000000000000000000000000 ;
        3510:  q   <=  32'b00000000000000000000000000000000 ;
        3511:  q   <=  32'b00000000000000000000000000000000 ;
        3512:  q   <=  32'b00000000000000000000000000000000 ;
        3513:  q   <=  32'b00000000000000000000000000000000 ;
        3514:  q   <=  32'b00000000000000000000000000000000 ;
        3515:  q   <=  32'b00000000000000000000000000000000 ;
        3516:  q   <=  32'b00000000000000000000000000000000 ;
        3517:  q   <=  32'b00000000000000000000000000000000 ;
        3518:  q   <=  32'b00000000000000000000000000000000 ;
        3519:  q   <=  32'b00000000000000000000000000000000 ;
        3520:  q   <=  32'b00000000000000000000000000000000 ;
        3521:  q   <=  32'b00000000000000000000000000000000 ;
        3522:  q   <=  32'b00000000000000000000000000000000 ;
        3523:  q   <=  32'b00000000000000000000000000000000 ;
        3524:  q   <=  32'b00000000000000000000000000000000 ;
        3525:  q   <=  32'b00000000000000000000000000000000 ;
        3526:  q   <=  32'b00000000000000000000000000000000 ;
        3527:  q   <=  32'b00000000000000000000000000000000 ;
        3528:  q   <=  32'b00000000000000000000000000000000 ;
        3529:  q   <=  32'b00000000000000000000000000000000 ;
        3530:  q   <=  32'b00000000000000000000000000000000 ;
        3531:  q   <=  32'b00000000000000000000000000000000 ;
        3532:  q   <=  32'b00000000000000000000000000000000 ;
        3533:  q   <=  32'b00000000000000000000000000000000 ;
        3534:  q   <=  32'b00000000000000000000000000000000 ;
        3535:  q   <=  32'b00000000000000000000000000000000 ;
        3536:  q   <=  32'b00000000000000000000000000000000 ;
        3537:  q   <=  32'b00000000000000000000000000000000 ;
        3538:  q   <=  32'b00000000000000000000000000000000 ;
        3539:  q   <=  32'b00000000000000000000000000000000 ;
        3540:  q   <=  32'b00000000000000000000000000000000 ;
        3541:  q   <=  32'b00000000000000000000000000000000 ;
        3542:  q   <=  32'b00000000000000000000000000000000 ;
        3543:  q   <=  32'b00000000000000000000000000000000 ;
        3544:  q   <=  32'b00000000000000000000000000000000 ;
        3545:  q   <=  32'b00000000000000000000000000000000 ;
        3546:  q   <=  32'b00000000000000000000000000000000 ;
        3547:  q   <=  32'b00000000000000000000000000000000 ;
        3548:  q   <=  32'b00000000000000000000000000000000 ;
        3549:  q   <=  32'b00000000000000000000000000000000 ;
        3550:  q   <=  32'b00000000000000000000000000000000 ;
        3551:  q   <=  32'b00000000000000000000000000000000 ;
        3552:  q   <=  32'b00111101101010000010000111100000 ;
        3553:  q   <=  32'b00111110100100010001100001110100 ;
        3554:  q   <=  32'b00111110111101111001001001001011 ;
        3555:  q   <=  32'b00111111001011101011101110100010 ;
        3556:  q   <=  32'b00111111011000010110010001010000 ;
        3557:  q   <=  32'b00111111100010011110000111101000 ;
        3558:  q   <=  32'b00111111101000101110110101100001 ;
        3559:  q   <=  32'b00111111101110111101010011100000 ;
        3560:  q   <=  32'b00111111110101001001100010110011 ;
        3561:  q   <=  32'b00111111111011010011100100100110 ;
        3562:  q   <=  32'b00111111111110100100100101111011 ;
        3563:  q   <=  32'b00111111111000011110111011100110 ;
        3564:  q   <=  32'b00111111110010011011011011010000 ;
        3565:  q   <=  32'b00111111101100011010000011110010 ;
        3566:  q   <=  32'b00111111100110011010110100000001 ;
        3567:  q   <=  32'b00111111100000011101101010110111 ;
        3568:  q   <=  32'b00111111010101000101001110011011 ;
        3569:  q   <=  32'b00111111001001010011001111111011 ;
        3570:  q   <=  32'b00111110111011001010110000001100 ;
        3571:  q   <=  32'b00111110100011110111001001100010 ;
        3572:  q   <=  32'b00111101110010101110011110101101 ;
        3573:  q   <=  32'b00000000000000000000000000000000 ;
        3574:  q   <=  32'b00000000000000000000000000000000 ;
        3575:  q   <=  32'b00000000000000000000000000000000 ;
        3576:  q   <=  32'b00000000000000000000000000000000 ;
        3577:  q   <=  32'b00000000000000000000000000000000 ;
        3578:  q   <=  32'b00000000000000000000000000000000 ;
        3579:  q   <=  32'b00000000000000000000000000000000 ;
        3580:  q   <=  32'b00000000000000000000000000000000 ;
        3581:  q   <=  32'b00000000000000000000000000000000 ;
        3582:  q   <=  32'b00000000000000000000000000000000 ;
        3583:  q   <=  32'b00000000000000000000000000000000 ;
        3584:  q   <=  32'b00000000000000000000000000000000 ;
        3585:  q   <=  32'b00000000000000000000000000000000 ;
        3586:  q   <=  32'b00000000000000000000000000000000 ;
        3587:  q   <=  32'b00000000000000000000000000000000 ;
        3588:  q   <=  32'b00000000000000000000000000000000 ;
        3589:  q   <=  32'b00000000000000000000000000000000 ;
        3590:  q   <=  32'b00000000000000000000000000000000 ;
        3591:  q   <=  32'b00000000000000000000000000000000 ;
        3592:  q   <=  32'b00000000000000000000000000000000 ;
        3593:  q   <=  32'b00000000000000000000000000000000 ;
        3594:  q   <=  32'b00000000000000000000000000000000 ;
        3595:  q   <=  32'b00000000000000000000000000000000 ;
        3596:  q   <=  32'b00000000000000000000000000000000 ;
        3597:  q   <=  32'b00000000000000000000000000000000 ;
        3598:  q   <=  32'b00000000000000000000000000000000 ;
        3599:  q   <=  32'b00000000000000000000000000000000 ;
        3600:  q   <=  32'b00000000000000000000000000000000 ;
        3601:  q   <=  32'b00000000000000000000000000000000 ;
        3602:  q   <=  32'b00000000000000000000000000000000 ;
        3603:  q   <=  32'b00000000000000000000000000000000 ;
        3604:  q   <=  32'b00000000000000000000000000000000 ;
        3605:  q   <=  32'b00000000000000000000000000000000 ;
        3606:  q   <=  32'b00000000000000000000000000000000 ;
        3607:  q   <=  32'b00000000000000000000000000000000 ;
        3608:  q   <=  32'b00000000000000000000000000000000 ;
        3609:  q   <=  32'b00000000000000000000000000000000 ;
        3610:  q   <=  32'b00000000000000000000000000000000 ;
        3611:  q   <=  32'b00000000000000000000000000000000 ;
        3612:  q   <=  32'b00000000000000000000000000000000 ;
        3613:  q   <=  32'b00000000000000000000000000000000 ;
        3614:  q   <=  32'b00000000000000000000000000000000 ;
        3615:  q   <=  32'b00000000000000000000000000000000 ;
        3616:  q   <=  32'b00000000000000000000000000000000 ;
        3617:  q   <=  32'b00000000000000000000000000000000 ;
        3618:  q   <=  32'b00000000000000000000000000000000 ;
        3619:  q   <=  32'b00000000000000000000000000000000 ;
        3620:  q   <=  32'b00000000000000000000000000000000 ;
        3621:  q   <=  32'b00000000000000000000000000000000 ;
        3622:  q   <=  32'b00000000000000000000000000000000 ;
        3623:  q   <=  32'b00000000000000000000000000000000 ;
        3624:  q   <=  32'b00000000000000000000000000000000 ;
        3625:  q   <=  32'b00000000000000000000000000000000 ;
        3626:  q   <=  32'b00000000000000000000000000000000 ;
        3627:  q   <=  32'b00000000000000000000000000000000 ;
        3628:  q   <=  32'b00000000000000000000000000000000 ;
        3629:  q   <=  32'b00000000000000000000000000000000 ;
        3630:  q   <=  32'b00000000000000000000000000000000 ;
        3631:  q   <=  32'b00000000000000000000000000000000 ;
        3632:  q   <=  32'b00000000000000000000000000000000 ;
        3633:  q   <=  32'b00000000000000000000000000000000 ;
        3634:  q   <=  32'b00000000000000000000000000000000 ;
        3635:  q   <=  32'b00000000000000000000000000000000 ;
        3636:  q   <=  32'b00000000000000000000000000000000 ;
        3637:  q   <=  32'b00000000000000000000000000000000 ;
        3638:  q   <=  32'b00000000000000000000000000000000 ;
        3639:  q   <=  32'b00000000000000000000000000000000 ;
        3640:  q   <=  32'b00000000000000000000000000000000 ;
        3641:  q   <=  32'b00000000000000000000000000000000 ;
        3642:  q   <=  32'b00000000000000000000000000000000 ;
        3643:  q   <=  32'b00000000000000000000000000000000 ;
        3644:  q   <=  32'b00000000000000000000000000000000 ;
        3645:  q   <=  32'b00000000000000000000000000000000 ;
        3646:  q   <=  32'b00000000000000000000000000000000 ;
        3647:  q   <=  32'b00000000000000000000000000000000 ;
        3648:  q   <=  32'b00000000000000000000000000000000 ;
        3649:  q   <=  32'b00000000000000000000000000000000 ;
        3650:  q   <=  32'b00000000000000000000000000000000 ;
        3651:  q   <=  32'b00000000000000000000000000000000 ;
        3652:  q   <=  32'b00000000000000000000000000000000 ;
        3653:  q   <=  32'b00000000000000000000000000000000 ;
        3654:  q   <=  32'b00000000000000000000000000000000 ;
        3655:  q   <=  32'b00000000000000000000000000000000 ;
        3656:  q   <=  32'b00000000000000000000000000000000 ;
        3657:  q   <=  32'b00000000000000000000000000000000 ;
        3658:  q   <=  32'b00000000000000000000000000000000 ;
        3659:  q   <=  32'b00000000000000000000000000000000 ;
        3660:  q   <=  32'b00000000000000000000000000000000 ;
        3661:  q   <=  32'b00000000000000000000000000000000 ;
        3662:  q   <=  32'b00000000000000000000000000000000 ;
        3663:  q   <=  32'b00000000000000000000000000000000 ;
        3664:  q   <=  32'b00000000000000000000000000000000 ;
        3665:  q   <=  32'b00000000000000000000000000000000 ;
        3666:  q   <=  32'b00000000000000000000000000000000 ;
        3667:  q   <=  32'b00000000000000000000000000000000 ;
        3668:  q   <=  32'b00000000000000000000000000000000 ;
        3669:  q   <=  32'b00000000000000000000000000000000 ;
        3670:  q   <=  32'b00000000000000000000000000000000 ;
        3671:  q   <=  32'b00000000000000000000000000000000 ;
        3672:  q   <=  32'b00000000000000000000000000000000 ;
        3673:  q   <=  32'b00000000000000000000000000000000 ;
        3674:  q   <=  32'b00000000000000000000000000000000 ;
        3675:  q   <=  32'b00000000000000000000000000000000 ;
        3676:  q   <=  32'b00000000000000000000000000000000 ;
        3677:  q   <=  32'b00000000000000000000000000000000 ;
        3678:  q   <=  32'b00000000000000000000000000000000 ;
        3679:  q   <=  32'b00000000000000000000000000000000 ;
        3680:  q   <=  32'b00000000000000000000000000000000 ;
        3681:  q   <=  32'b00000000000000000000000000000000 ;
        3682:  q   <=  32'b00000000000000000000000000000000 ;
        3683:  q   <=  32'b00000000000000000000000000000000 ;
        3684:  q   <=  32'b00000000000000000000000000000000 ;
        3685:  q   <=  32'b00000000000000000000000000000000 ;
        3686:  q   <=  32'b00000000000000000000000000000000 ;
        3687:  q   <=  32'b00000000000000000000000000000000 ;
        3688:  q   <=  32'b00000000000000000000000000000000 ;
        3689:  q   <=  32'b00000000000000000000000000000000 ;
        3690:  q   <=  32'b00000000000000000000000000000000 ;
        3691:  q   <=  32'b00000000000000000000000000000000 ;
        3692:  q   <=  32'b00000000000000000000000000000000 ;
        3693:  q   <=  32'b00000000000000000000000000000000 ;
        3694:  q   <=  32'b00000000000000000000000000000000 ;
        3695:  q   <=  32'b00000000000000000000000000000000 ;
        3696:  q   <=  32'b00000000000000000000000000000000 ;
        3697:  q   <=  32'b00000000000000000000000000000000 ;
        3698:  q   <=  32'b00000000000000000000000000000000 ;
        3699:  q   <=  32'b00000000000000000000000000000000 ;
        3700:  q   <=  32'b00000000000000000000000000000000 ;
        3701:  q   <=  32'b00000000000000000000000000000000 ;
        3702:  q   <=  32'b00000000000000000000000000000000 ;
        3703:  q   <=  32'b00000000000000000000000000000000 ;
        3704:  q   <=  32'b00000000000000000000000000000000 ;
        3705:  q   <=  32'b00000000000000000000000000000000 ;
        3706:  q   <=  32'b00000000000000000000000000000000 ;
        3707:  q   <=  32'b00000000000000000000000000000000 ;
        3708:  q   <=  32'b00000000000000000000000000000000 ;
        3709:  q   <=  32'b00000000000000000000000000000000 ;
        3710:  q   <=  32'b00000000000000000000000000000000 ;
        3711:  q   <=  32'b00000000000000000000000000000000 ;
        3712:  q   <=  32'b00000000000000000000000000000000 ;
        3713:  q   <=  32'b00000000000000000000000000000000 ;
        3714:  q   <=  32'b00000000000000000000000000000000 ;
        3715:  q   <=  32'b00000000000000000000000000000000 ;
        3716:  q   <=  32'b00000000000000000000000000000000 ;
        3717:  q   <=  32'b00000000000000000000000000000000 ;
        3718:  q   <=  32'b00000000000000000000000000000000 ;
        3719:  q   <=  32'b00000000000000000000000000000000 ;
        3720:  q   <=  32'b00000000000000000000000000000000 ;
        3721:  q   <=  32'b00000000000000000000000000000000 ;
        3722:  q   <=  32'b00000000000000000000000000000000 ;
        3723:  q   <=  32'b00000000000000000000000000000000 ;
        3724:  q   <=  32'b00000000000000000000000000000000 ;
        3725:  q   <=  32'b00000000000000000000000000000000 ;
        3726:  q   <=  32'b00000000000000000000000000000000 ;
        3727:  q   <=  32'b00000000000000000000000000000000 ;
        3728:  q   <=  32'b00000000000000000000000000000000 ;
        3729:  q   <=  32'b00000000000000000000000000000000 ;
        3730:  q   <=  32'b00000000000000000000000000000000 ;
        3731:  q   <=  32'b00000000000000000000000000000000 ;
        3732:  q   <=  32'b00000000000000000000000000000000 ;
        3733:  q   <=  32'b00000000000000000000000000000000 ;
        3734:  q   <=  32'b00000000000000000000000000000000 ;
        3735:  q   <=  32'b00000000000000000000000000000000 ;
        3736:  q   <=  32'b00000000000000000000000000000000 ;
        3737:  q   <=  32'b00000000000000000000000000000000 ;
        3738:  q   <=  32'b00000000000000000000000000000000 ;
        3739:  q   <=  32'b00000000000000000000000000000000 ;
        3740:  q   <=  32'b00000000000000000000000000000000 ;
        3741:  q   <=  32'b00000000000000000000000000000000 ;
        3742:  q   <=  32'b00000000000000000000000000000000 ;
        3743:  q   <=  32'b00000000000000000000000000000000 ;
        3744:  q   <=  32'b00000000000000000000000000000000 ;
        3745:  q   <=  32'b00000000000000000000000000000000 ;
        3746:  q   <=  32'b00000000000000000000000000000000 ;
        3747:  q   <=  32'b00000000000000000000000000000000 ;
        3748:  q   <=  32'b00000000000000000000000000000000 ;
        3749:  q   <=  32'b00000000000000000000000000000000 ;
        3750:  q   <=  32'b00000000000000000000000000000000 ;
        3751:  q   <=  32'b00000000000000000000000000000000 ;
        3752:  q   <=  32'b00000000000000000000000000000000 ;
        3753:  q   <=  32'b00000000000000000000000000000000 ;
        3754:  q   <=  32'b00000000000000000000000000000000 ;
        3755:  q   <=  32'b00000000000000000000000000000000 ;
        3756:  q   <=  32'b00000000000000000000000000000000 ;
        3757:  q   <=  32'b00000000000000000000000000000000 ;
        3758:  q   <=  32'b00000000000000000000000000000000 ;
        3759:  q   <=  32'b00000000000000000000000000000000 ;
        3760:  q   <=  32'b00000000000000000000000000000000 ;
        3761:  q   <=  32'b00000000000000000000000000000000 ;
        3762:  q   <=  32'b00000000000000000000000000000000 ;
        3763:  q   <=  32'b00000000000000000000000000000000 ;
        3764:  q   <=  32'b00000000000000000000000000000000 ;
        3765:  q   <=  32'b00000000000000000000000000000000 ;
        3766:  q   <=  32'b00000000000000000000000000000000 ;
        3767:  q   <=  32'b00000000000000000000000000000000 ;
        3768:  q   <=  32'b00000000000000000000000000000000 ;
        3769:  q   <=  32'b00000000000000000000000000000000 ;
        3770:  q   <=  32'b00000000000000000000000000000000 ;
        3771:  q   <=  32'b00000000000000000000000000000000 ;
        3772:  q   <=  32'b00000000000000000000000000000000 ;
        3773:  q   <=  32'b00000000000000000000000000000000 ;
        3774:  q   <=  32'b00000000000000000000000000000000 ;
        3775:  q   <=  32'b00000000000000000000000000000000 ;
        3776:  q   <=  32'b00000000000000000000000000000000 ;
        3777:  q   <=  32'b00000000000000000000000000000000 ;
        3778:  q   <=  32'b00000000000000000000000000000000 ;
        3779:  q   <=  32'b00000000000000000000000000000000 ;
        3780:  q   <=  32'b00000000000000000000000000000000 ;
        3781:  q   <=  32'b00000000000000000000000000000000 ;
        3782:  q   <=  32'b00000000000000000000000000000000 ;
        3783:  q   <=  32'b00000000000000000000000000000000 ;
        3784:  q   <=  32'b00000000000000000000000000000000 ;
        3785:  q   <=  32'b00000000000000000000000000000000 ;
        3786:  q   <=  32'b00000000000000000000000000000000 ;
        3787:  q   <=  32'b00000000000000000000000000000000 ;
        3788:  q   <=  32'b00000000000000000000000000000000 ;
        3789:  q   <=  32'b00000000000000000000000000000000 ;
        3790:  q   <=  32'b00000000000000000000000000000000 ;
        3791:  q   <=  32'b00000000000000000000000000000000 ;
        3792:  q   <=  32'b00000000000000000000000000000000 ;
        3793:  q   <=  32'b00000000000000000000000000000000 ;
        3794:  q   <=  32'b00000000000000000000000000000000 ;
        3795:  q   <=  32'b00000000000000000000000000000000 ;
        3796:  q   <=  32'b00000000000000000000000000000000 ;
        3797:  q   <=  32'b00000000000000000000000000000000 ;
        3798:  q   <=  32'b00000000000000000000000000000000 ;
        3799:  q   <=  32'b00000000000000000000000000000000 ;
        3800:  q   <=  32'b00000000000000000000000000000000 ;
        3801:  q   <=  32'b00000000000000000000000000000000 ;
        3802:  q   <=  32'b00000000000000000000000000000000 ;
        3803:  q   <=  32'b00000000000000000000000000000000 ;
        3804:  q   <=  32'b00000000000000000000000000000000 ;
        3805:  q   <=  32'b00000000000000000000000000000000 ;
        3806:  q   <=  32'b00000000000000000000000000000000 ;
        3807:  q   <=  32'b00000000000000000000000000000000 ;
        3808:  q   <=  32'b00000000000000000000000000000000 ;
        3809:  q   <=  32'b00000000000000000000000000000000 ;
        3810:  q   <=  32'b00000000000000000000000000000000 ;
        3811:  q   <=  32'b00000000000000000000000000000000 ;
        3812:  q   <=  32'b00000000000000000000000000000000 ;
        3813:  q   <=  32'b00000000000000000000000000000000 ;
        3814:  q   <=  32'b00000000000000000000000000000000 ;
        3815:  q   <=  32'b00000000000000000000000000000000 ;
        3816:  q   <=  32'b00000000000000000000000000000000 ;
        3817:  q   <=  32'b00000000000000000000000000000000 ;
        3818:  q   <=  32'b00111101001101101101000010010100 ;
        3819:  q   <=  32'b00111110011100001000100011001101 ;
        3820:  q   <=  32'b00111110110110010010010010111100 ;
        3821:  q   <=  32'b00111111000111001011111000011011 ;
        3822:  q   <=  32'b00111111010011001010010111111100 ;
        3823:  q   <=  32'b00111111011111000100101010010000 ;
        3824:  q   <=  32'b00111111100101011101011000110010 ;
        3825:  q   <=  32'b00111111101011010110011000000010 ;
        3826:  q   <=  32'b00111111110001001101010011111100 ;
        3827:  q   <=  32'b00111111110111000010001101100111 ;
        3828:  q   <=  32'b00111111111100110101000110000101 ;
        3829:  q   <=  32'b00111111111101011010000001100110 ;
        3830:  q   <=  32'b00111111110111101011001000011010 ;
        3831:  q   <=  32'b00111111110001111110001101010100 ;
        3832:  q   <=  32'b00111111101100010011001111010010 ;
        3833:  q   <=  32'b00111111100110101010001101010110 ;
        3834:  q   <=  32'b00111111100001000011000110011111 ;
        3835:  q   <=  32'b00111111010110111011110011100000 ;
        3836:  q   <=  32'b00111111001011110101001100010010 ;
        3837:  q   <=  32'b00111111000000110010010101011010 ;
        3838:  q   <=  32'b00111110101011100110011001111110 ;
        3839:  q   <=  32'b00111110001011011111000100100011 ;
        3840:  q   <=  32'b00000000000000000000000000000000 ;
        3841:  q   <=  32'b00000000000000000000000000000000 ;
        3842:  q   <=  32'b00000000000000000000000000000000 ;
        3843:  q   <=  32'b00000000000000000000000000000000 ;
        3844:  q   <=  32'b00000000000000000000000000000000 ;
        3845:  q   <=  32'b00000000000000000000000000000000 ;
        3846:  q   <=  32'b00000000000000000000000000000000 ;
        3847:  q   <=  32'b00000000000000000000000000000000 ;
        3848:  q   <=  32'b00000000000000000000000000000000 ;
        3849:  q   <=  32'b00000000000000000000000000000000 ;
        3850:  q   <=  32'b00000000000000000000000000000000 ;
        3851:  q   <=  32'b00000000000000000000000000000000 ;
        3852:  q   <=  32'b00000000000000000000000000000000 ;
        3853:  q   <=  32'b00000000000000000000000000000000 ;
        3854:  q   <=  32'b00000000000000000000000000000000 ;
        3855:  q   <=  32'b00000000000000000000000000000000 ;
        3856:  q   <=  32'b00000000000000000000000000000000 ;
        3857:  q   <=  32'b00000000000000000000000000000000 ;
        3858:  q   <=  32'b00000000000000000000000000000000 ;
        3859:  q   <=  32'b00000000000000000000000000000000 ;
        3860:  q   <=  32'b00000000000000000000000000000000 ;
        3861:  q   <=  32'b00000000000000000000000000000000 ;
        3862:  q   <=  32'b00000000000000000000000000000000 ;
        3863:  q   <=  32'b00000000000000000000000000000000 ;
        3864:  q   <=  32'b00000000000000000000000000000000 ;
        3865:  q   <=  32'b00000000000000000000000000000000 ;
        3866:  q   <=  32'b00000000000000000000000000000000 ;
        3867:  q   <=  32'b00000000000000000000000000000000 ;
        3868:  q   <=  32'b00000000000000000000000000000000 ;
        3869:  q   <=  32'b00000000000000000000000000000000 ;
        3870:  q   <=  32'b00000000000000000000000000000000 ;
        3871:  q   <=  32'b00000000000000000000000000000000 ;
        3872:  q   <=  32'b00000000000000000000000000000000 ;
        3873:  q   <=  32'b00000000000000000000000000000000 ;
        3874:  q   <=  32'b00000000000000000000000000000000 ;
        3875:  q   <=  32'b00000000000000000000000000000000 ;
        3876:  q   <=  32'b00000000000000000000000000000000 ;
        3877:  q   <=  32'b00000000000000000000000000000000 ;
        3878:  q   <=  32'b00000000000000000000000000000000 ;
        3879:  q   <=  32'b00000000000000000000000000000000 ;
        3880:  q   <=  32'b00000000000000000000000000000000 ;
        3881:  q   <=  32'b00000000000000000000000000000000 ;
        3882:  q   <=  32'b00000000000000000000000000000000 ;
        3883:  q   <=  32'b00000000000000000000000000000000 ;
        3884:  q   <=  32'b00000000000000000000000000000000 ;
        3885:  q   <=  32'b00000000000000000000000000000000 ;
        3886:  q   <=  32'b00000000000000000000000000000000 ;
        3887:  q   <=  32'b00000000000000000000000000000000 ;
        3888:  q   <=  32'b00000000000000000000000000000000 ;
        3889:  q   <=  32'b00000000000000000000000000000000 ;
        3890:  q   <=  32'b00000000000000000000000000000000 ;
        3891:  q   <=  32'b00000000000000000000000000000000 ;
        3892:  q   <=  32'b00000000000000000000000000000000 ;
        3893:  q   <=  32'b00000000000000000000000000000000 ;
        3894:  q   <=  32'b00000000000000000000000000000000 ;
        3895:  q   <=  32'b00000000000000000000000000000000 ;
        3896:  q   <=  32'b00000000000000000000000000000000 ;
        3897:  q   <=  32'b00000000000000000000000000000000 ;
        3898:  q   <=  32'b00000000000000000000000000000000 ;
        3899:  q   <=  32'b00000000000000000000000000000000 ;
        3900:  q   <=  32'b00000000000000000000000000000000 ;
        3901:  q   <=  32'b00000000000000000000000000000000 ;
        3902:  q   <=  32'b00000000000000000000000000000000 ;
        3903:  q   <=  32'b00000000000000000000000000000000 ;
        3904:  q   <=  32'b00000000000000000000000000000000 ;
        3905:  q   <=  32'b00000000000000000000000000000000 ;
        3906:  q   <=  32'b00000000000000000000000000000000 ;
        3907:  q   <=  32'b00000000000000000000000000000000 ;
        3908:  q   <=  32'b00000000000000000000000000000000 ;
        3909:  q   <=  32'b00000000000000000000000000000000 ;
        3910:  q   <=  32'b00000000000000000000000000000000 ;
        3911:  q   <=  32'b00000000000000000000000000000000 ;
        3912:  q   <=  32'b00000000000000000000000000000000 ;
        3913:  q   <=  32'b00000000000000000000000000000000 ;
        3914:  q   <=  32'b00000000000000000000000000000000 ;
        3915:  q   <=  32'b00000000000000000000000000000000 ;
        3916:  q   <=  32'b00000000000000000000000000000000 ;
        3917:  q   <=  32'b00000000000000000000000000000000 ;
        3918:  q   <=  32'b00000000000000000000000000000000 ;
        3919:  q   <=  32'b00000000000000000000000000000000 ;
        3920:  q   <=  32'b00000000000000000000000000000000 ;
        3921:  q   <=  32'b00000000000000000000000000000000 ;
        3922:  q   <=  32'b00000000000000000000000000000000 ;
        3923:  q   <=  32'b00000000000000000000000000000000 ;
        3924:  q   <=  32'b00000000000000000000000000000000 ;
        3925:  q   <=  32'b00000000000000000000000000000000 ;
        3926:  q   <=  32'b00000000000000000000000000000000 ;
        3927:  q   <=  32'b00000000000000000000000000000000 ;
        3928:  q   <=  32'b00000000000000000000000000000000 ;
        3929:  q   <=  32'b00000000000000000000000000000000 ;
        3930:  q   <=  32'b00000000000000000000000000000000 ;
        3931:  q   <=  32'b00000000000000000000000000000000 ;
        3932:  q   <=  32'b00000000000000000000000000000000 ;
        3933:  q   <=  32'b00000000000000000000000000000000 ;
        3934:  q   <=  32'b00000000000000000000000000000000 ;
        3935:  q   <=  32'b00000000000000000000000000000000 ;
        3936:  q   <=  32'b00000000000000000000000000000000 ;
        3937:  q   <=  32'b00000000000000000000000000000000 ;
        3938:  q   <=  32'b00000000000000000000000000000000 ;
        3939:  q   <=  32'b00000000000000000000000000000000 ;
        3940:  q   <=  32'b00000000000000000000000000000000 ;
        3941:  q   <=  32'b00000000000000000000000000000000 ;
        3942:  q   <=  32'b00000000000000000000000000000000 ;
        3943:  q   <=  32'b00000000000000000000000000000000 ;
        3944:  q   <=  32'b00000000000000000000000000000000 ;
        3945:  q   <=  32'b00000000000000000000000000000000 ;
        3946:  q   <=  32'b00000000000000000000000000000000 ;
        3947:  q   <=  32'b00000000000000000000000000000000 ;
        3948:  q   <=  32'b00000000000000000000000000000000 ;
        3949:  q   <=  32'b00000000000000000000000000000000 ;
        3950:  q   <=  32'b00000000000000000000000000000000 ;
        3951:  q   <=  32'b00000000000000000000000000000000 ;
        3952:  q   <=  32'b00000000000000000000000000000000 ;
        3953:  q   <=  32'b00000000000000000000000000000000 ;
        3954:  q   <=  32'b00000000000000000000000000000000 ;
        3955:  q   <=  32'b00000000000000000000000000000000 ;
        3956:  q   <=  32'b00000000000000000000000000000000 ;
        3957:  q   <=  32'b00000000000000000000000000000000 ;
        3958:  q   <=  32'b00000000000000000000000000000000 ;
        3959:  q   <=  32'b00000000000000000000000000000000 ;
        3960:  q   <=  32'b00000000000000000000000000000000 ;
        3961:  q   <=  32'b00000000000000000000000000000000 ;
        3962:  q   <=  32'b00000000000000000000000000000000 ;
        3963:  q   <=  32'b00000000000000000000000000000000 ;
        3964:  q   <=  32'b00000000000000000000000000000000 ;
        3965:  q   <=  32'b00000000000000000000000000000000 ;
        3966:  q   <=  32'b00000000000000000000000000000000 ;
        3967:  q   <=  32'b00000000000000000000000000000000 ;
        3968:  q   <=  32'b00000000000000000000000000000000 ;
        3969:  q   <=  32'b00000000000000000000000000000000 ;
        3970:  q   <=  32'b00000000000000000000000000000000 ;
        3971:  q   <=  32'b00000000000000000000000000000000 ;
        3972:  q   <=  32'b00000000000000000000000000000000 ;
        3973:  q   <=  32'b00000000000000000000000000000000 ;
        3974:  q   <=  32'b00000000000000000000000000000000 ;
        3975:  q   <=  32'b00000000000000000000000000000000 ;
        3976:  q   <=  32'b00000000000000000000000000000000 ;
        3977:  q   <=  32'b00000000000000000000000000000000 ;
        3978:  q   <=  32'b00000000000000000000000000000000 ;
        3979:  q   <=  32'b00000000000000000000000000000000 ;
        3980:  q   <=  32'b00000000000000000000000000000000 ;
        3981:  q   <=  32'b00000000000000000000000000000000 ;
        3982:  q   <=  32'b00000000000000000000000000000000 ;
        3983:  q   <=  32'b00000000000000000000000000000000 ;
        3984:  q   <=  32'b00000000000000000000000000000000 ;
        3985:  q   <=  32'b00000000000000000000000000000000 ;
        3986:  q   <=  32'b00000000000000000000000000000000 ;
        3987:  q   <=  32'b00000000000000000000000000000000 ;
        3988:  q   <=  32'b00000000000000000000000000000000 ;
        3989:  q   <=  32'b00000000000000000000000000000000 ;
        3990:  q   <=  32'b00000000000000000000000000000000 ;
        3991:  q   <=  32'b00000000000000000000000000000000 ;
        3992:  q   <=  32'b00000000000000000000000000000000 ;
        3993:  q   <=  32'b00000000000000000000000000000000 ;
        3994:  q   <=  32'b00000000000000000000000000000000 ;
        3995:  q   <=  32'b00000000000000000000000000000000 ;
        3996:  q   <=  32'b00000000000000000000000000000000 ;
        3997:  q   <=  32'b00000000000000000000000000000000 ;
        3998:  q   <=  32'b00000000000000000000000000000000 ;
        3999:  q   <=  32'b00000000000000000000000000000000 ;
        4000:  q   <=  32'b00000000000000000000000000000000 ;
        4001:  q   <=  32'b00000000000000000000000000000000 ;
        4002:  q   <=  32'b00000000000000000000000000000000 ;
        4003:  q   <=  32'b00000000000000000000000000000000 ;
        4004:  q   <=  32'b00000000000000000000000000000000 ;
        4005:  q   <=  32'b00000000000000000000000000000000 ;
        4006:  q   <=  32'b00000000000000000000000000000000 ;
        4007:  q   <=  32'b00000000000000000000000000000000 ;
        4008:  q   <=  32'b00000000000000000000000000000000 ;
        4009:  q   <=  32'b00000000000000000000000000000000 ;
        4010:  q   <=  32'b00000000000000000000000000000000 ;
        4011:  q   <=  32'b00000000000000000000000000000000 ;
        4012:  q   <=  32'b00000000000000000000000000000000 ;
        4013:  q   <=  32'b00000000000000000000000000000000 ;
        4014:  q   <=  32'b00000000000000000000000000000000 ;
        4015:  q   <=  32'b00000000000000000000000000000000 ;
        4016:  q   <=  32'b00000000000000000000000000000000 ;
        4017:  q   <=  32'b00000000000000000000000000000000 ;
        4018:  q   <=  32'b00000000000000000000000000000000 ;
        4019:  q   <=  32'b00000000000000000000000000000000 ;
        4020:  q   <=  32'b00000000000000000000000000000000 ;
        4021:  q   <=  32'b00000000000000000000000000000000 ;
        4022:  q   <=  32'b00000000000000000000000000000000 ;
        4023:  q   <=  32'b00000000000000000000000000000000 ;
        4024:  q   <=  32'b00000000000000000000000000000000 ;
        4025:  q   <=  32'b00000000000000000000000000000000 ;
        4026:  q   <=  32'b00000000000000000000000000000000 ;
        4027:  q   <=  32'b00000000000000000000000000000000 ;
        4028:  q   <=  32'b00000000000000000000000000000000 ;
        4029:  q   <=  32'b00000000000000000000000000000000 ;
        4030:  q   <=  32'b00000000000000000000000000000000 ;
        4031:  q   <=  32'b00000000000000000000000000000000 ;
        4032:  q   <=  32'b00000000000000000000000000000000 ;
        4033:  q   <=  32'b00000000000000000000000000000000 ;
        4034:  q   <=  32'b00000000000000000000000000000000 ;
        4035:  q   <=  32'b00000000000000000000000000000000 ;
        4036:  q   <=  32'b00000000000000000000000000000000 ;
        4037:  q   <=  32'b00000000000000000000000000000000 ;
        4038:  q   <=  32'b00000000000000000000000000000000 ;
        4039:  q   <=  32'b00000000000000000000000000000000 ;
        4040:  q   <=  32'b00000000000000000000000000000000 ;
        4041:  q   <=  32'b00000000000000000000000000000000 ;
        4042:  q   <=  32'b00000000000000000000000000000000 ;
        4043:  q   <=  32'b00000000000000000000000000000000 ;
        4044:  q   <=  32'b00000000000000000000000000000000 ;
        4045:  q   <=  32'b00000000000000000000000000000000 ;
        4046:  q   <=  32'b00000000000000000000000000000000 ;
        4047:  q   <=  32'b00000000000000000000000000000000 ;
        4048:  q   <=  32'b00000000000000000000000000000000 ;
        4049:  q   <=  32'b00000000000000000000000000000000 ;
        4050:  q   <=  32'b00000000000000000000000000000000 ;
        4051:  q   <=  32'b00000000000000000000000000000000 ;
        4052:  q   <=  32'b00000000000000000000000000000000 ;
        4053:  q   <=  32'b00000000000000000000000000000000 ;
        4054:  q   <=  32'b00000000000000000000000000000000 ;
        4055:  q   <=  32'b00000000000000000000000000000000 ;
        4056:  q   <=  32'b00000000000000000000000000000000 ;
        4057:  q   <=  32'b00000000000000000000000000000000 ;
        4058:  q   <=  32'b00000000000000000000000000000000 ;
        4059:  q   <=  32'b00000000000000000000000000000000 ;
        4060:  q   <=  32'b00000000000000000000000000000000 ;
        4061:  q   <=  32'b00000000000000000000000000000000 ;
        4062:  q   <=  32'b00000000000000000000000000000000 ;
        4063:  q   <=  32'b00000000000000000000000000000000 ;
        4064:  q   <=  32'b00000000000000000000000000000000 ;
        4065:  q   <=  32'b00000000000000000000000000000000 ;
        4066:  q   <=  32'b00000000000000000000000000000000 ;
        4067:  q   <=  32'b00000000000000000000000000000000 ;
        4068:  q   <=  32'b00000000000000000000000000000000 ;
        4069:  q   <=  32'b00000000000000000000000000000000 ;
        4070:  q   <=  32'b00000000000000000000000000000000 ;
        4071:  q   <=  32'b00000000000000000000000000000000 ;
        4072:  q   <=  32'b00000000000000000000000000000000 ;
        4073:  q   <=  32'b00000000000000000000000000000000 ;
        4074:  q   <=  32'b00000000000000000000000000000000 ;
        4075:  q   <=  32'b00000000000000000000000000000000 ;
        4076:  q   <=  32'b00000000000000000000000000000000 ;
        4077:  q   <=  32'b00000000000000000000000000000000 ;
        4078:  q   <=  32'b00000000000000000000000000000000 ;
        4079:  q   <=  32'b00000000000000000000000000000000 ;
        4080:  q   <=  32'b00000000000000000000000000000000 ;
        4081:  q   <=  32'b00000000000000000000000000000000 ;
        4082:  q   <=  32'b00000000000000000000000000000000 ;
        4083:  q   <=  32'b00000000000000000000000000000000 ;
        4084:  q   <=  32'b00000000000000000000000000000000 ;
        4085:  q   <=  32'b00000000000000000000000000000000 ;
        4086:  q   <=  32'b00000000000000000000000000000000 ;
        4087:  q   <=  32'b00000000000000000000000000000000 ;
        4088:  q   <=  32'b00000000000000000000000000000000 ;
        4089:  q   <=  32'b00000000000000000000000000000000 ;
        4090:  q   <=  32'b00000000000000000000000000000000 ;
        4091:  q   <=  32'b00000000000000000000000000000000 ;
        4092:  q   <=  32'b00000000000000000000000000000000 ;
        4093:  q   <=  32'b00000000000000000000000000000000 ;
        4094:  q   <=  32'b00000000000000000000000000000000 ;
        4095:  q   <=  32'b00000000000000000000000000000000;
        default: q <= 0;
    endcase
end
endmodule
