module mem_mantissa (clk, addr, cen, wen, data, q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;// Note
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00111000110111100101010011100110 ;
        2:  q   <=  32'b00111001010111100100110111110100 ;
        3:  q   <=  32'b00111001101001101011010101000001 ;
        4:  q   <=  32'b00111001110111100100000000010001 ;
        5:  q   <=  32'b00111010000010101110001110110100 ;
        6:  q   <=  32'b00111010001001101010010110100101 ;
        7:  q   <=  32'b00111010010000100110010111011010 ;
        8:  q   <=  32'b00111010010111100010010001010100 ;
        9:  q   <=  32'b00111010011110011110000100010011 ;
        10:  q   <=  32'b00111010100010101100111000001011 ;
        11:  q   <=  32'b00111010100110001010101010110000 ;
        12:  q   <=  32'b00111010101001101000011001110111 ;
        13:  q   <=  32'b00111010101101000110000101100010 ;
        14:  q   <=  32'b00111010110000100011101101101111 ;
        15:  q   <=  32'b00111010110100000001010010100000 ;
        16:  q   <=  32'b00111010110111011110110011110100 ;
        17:  q   <=  32'b00111010111010111100010001101011 ;
        18:  q   <=  32'b00111010111110011001101100000110 ;
        19:  q   <=  32'b00111011000000111011100001100010 ;
        20:  q   <=  32'b00111011000010101010001011010011 ;
        21:  q   <=  32'b00111011000100011000110011010110 ;
        22:  q   <=  32'b00111011000110000111011001101011 ;
        23:  q   <=  32'b00111011000111110101111110010010 ;
        24:  q   <=  32'b00111011001001100100100001001011 ;
        25:  q   <=  32'b00111011001011010011000010010110 ;
        26:  q   <=  32'b00111011001101000001100001110011 ;
        27:  q   <=  32'b00111011001110101111111111100011 ;
        28:  q   <=  32'b00111011010000011110011011100100 ;
        29:  q   <=  32'b00111011010010001100110101111000 ;
        30:  q   <=  32'b00111011010011111011001110011111 ;
        31:  q   <=  32'b00111011010101101001100101011000 ;
        32:  q   <=  32'b00111011010111010111111010100011 ;
        33:  q   <=  32'b00111011011001000110001110000001 ;
        34:  q   <=  32'b00111011011010110100011111110001 ;
        35:  q   <=  32'b00111011011100100010101111110101 ;
        36:  q   <=  32'b00111011011110010000111110001010 ;
        37:  q   <=  32'b00111011011111111111001010110011 ;
        38:  q   <=  32'b00111011100000110110101010110111 ;
        39:  q   <=  32'b00111011100001101101101111011110 ;
        40:  q   <=  32'b00111011100010100100110011001111 ;
        41:  q   <=  32'b00111011100011011011110110001001 ;
        42:  q   <=  32'b00111011100100010010111000001100 ;
        43:  q   <=  32'b00111011100101001001111001011001 ;
        44:  q   <=  32'b00111011100110000000111001110000 ;
        45:  q   <=  32'b00111011100110110111111001010000 ;
        46:  q   <=  32'b00111011100111101110110111111010 ;
        47:  q   <=  32'b00111011101000100101110101101101 ;
        48:  q   <=  32'b00111011101001011100110010101011 ;
        49:  q   <=  32'b00111011101010010011101110110001 ;
        50:  q   <=  32'b00111011101011001010101010000010 ;
        51:  q   <=  32'b00111011101100000001100100011100 ;
        52:  q   <=  32'b00111011101100111000011110000000 ;
        53:  q   <=  32'b00111011101101101111010110101110 ;
        54:  q   <=  32'b00111011101110100110001110100110 ;
        55:  q   <=  32'b00111011101111011101000101100111 ;
        56:  q   <=  32'b00111011110000010011111011110011 ;
        57:  q   <=  32'b00111011110001001010110001001000 ;
        58:  q   <=  32'b00111011110010000001100101100111 ;
        59:  q   <=  32'b00111011110010111000011001010001 ;
        60:  q   <=  32'b00111011110011101111001100000100 ;
        61:  q   <=  32'b00111011110100100101111110000001 ;
        62:  q   <=  32'b00111011110101011100101111001000 ;
        63:  q   <=  32'b00111011110110010011011111011001 ;
        64:  q   <=  32'b00111011110111001010001110110101 ;
        65:  q   <=  32'b00111011111000000000111101011010 ;
        66:  q   <=  32'b00111011111000110111101011001010 ;
        67:  q   <=  32'b00111011111001101110011000000011 ;
        68:  q   <=  32'b00111011111010100101000100000111 ;
        69:  q   <=  32'b00111011111011011011101111010101 ;
        70:  q   <=  32'b00111011111100010010011001101110 ;
        71:  q   <=  32'b00111011111101001001000011010000 ;
        72:  q   <=  32'b00111011111101111111101011111101 ;
        73:  q   <=  32'b00111011111110110110010011110101 ;
        74:  q   <=  32'b00111011111111101100111010110110 ;
        75:  q   <=  32'b00111100000000010001110000100001 ;
        76:  q   <=  32'b00111100000000101101000011001100 ;
        77:  q   <=  32'b00111100000001001000010101011100 ;
        78:  q   <=  32'b00111100000001100011100111010010 ;
        79:  q   <=  32'b00111100000001111110111000101101 ;
        80:  q   <=  32'b00111100000010011010001001101101 ;
        81:  q   <=  32'b00111100000010110101011010010010 ;
        82:  q   <=  32'b00111100000011010000101010011101 ;
        83:  q   <=  32'b00111100000011101011111010001101 ;
        84:  q   <=  32'b00111100000100000111001001100010 ;
        85:  q   <=  32'b00111100000100100010011000011100 ;
        86:  q   <=  32'b00111100000100111101100110111100 ;
        87:  q   <=  32'b00111100000101011000110101000001 ;
        88:  q   <=  32'b00111100000101110100000010101100 ;
        89:  q   <=  32'b00111100000110001111001111111100 ;
        90:  q   <=  32'b00111100000110101010011100110001 ;
        91:  q   <=  32'b00111100000111000101101001001100 ;
        92:  q   <=  32'b00111100000111100000110101001100 ;
        93:  q   <=  32'b00111100000111111100000000110001 ;
        94:  q   <=  32'b00111100001000010111001011111100 ;
        95:  q   <=  32'b00111100001000110010010110101100 ;
        96:  q   <=  32'b00111100001001001101100001000010 ;
        97:  q   <=  32'b00111100001001101000101010111101 ;
        98:  q   <=  32'b00111100001010000011110100011110 ;
        99:  q   <=  32'b00111100001010011110111101100100 ;
        100:  q   <=  32'b00111100001010111010000110010000 ;
        101:  q   <=  32'b00111100001011010101001110100001 ;
        102:  q   <=  32'b00111100001011110000010110011000 ;
        103:  q   <=  32'b00111100001100001011011101110100 ;
        104:  q   <=  32'b00111100001100100110100100110110 ;
        105:  q   <=  32'b00111100001101000001101011011101 ;
        106:  q   <=  32'b00111100001101011100110001101010 ;
        107:  q   <=  32'b00111100001101110111110111011101 ;
        108:  q   <=  32'b00111100001110010010111100110101 ;
        109:  q   <=  32'b00111100001110101110000001110011 ;
        110:  q   <=  32'b00111100001111001001000110010110 ;
        111:  q   <=  32'b00111100001111100100001010011111 ;
        112:  q   <=  32'b00111100001111111111001110001110 ;
        113:  q   <=  32'b00111100010000011010010001100010 ;
        114:  q   <=  32'b00111100010000110101010100011100 ;
        115:  q   <=  32'b00111100010001010000010110111100 ;
        116:  q   <=  32'b00111100010001101011011001000001 ;
        117:  q   <=  32'b00111100010010000110011010101101 ;
        118:  q   <=  32'b00111100010010100001011011111101 ;
        119:  q   <=  32'b00111100010010111100011100110100 ;
        120:  q   <=  32'b00111100010011010111011101010000 ;
        121:  q   <=  32'b00111100010011110010011101010011 ;
        122:  q   <=  32'b00111100010100001101011100111010 ;
        123:  q   <=  32'b00111100010100101000011100001000 ;
        124:  q   <=  32'b00111100010101000011011010111100 ;
        125:  q   <=  32'b00111100010101011110011001010101 ;
        126:  q   <=  32'b00111100010101111001010111010100 ;
        127:  q   <=  32'b00111100010110010100010100111001 ;
        128:  q   <=  32'b00111100010110101111010010000100 ;
        129:  q   <=  32'b00111100010111001010001110110101 ;
        130:  q   <=  32'b00111100010111100101001011001011 ;
        131:  q   <=  32'b00111100011000000000000111001000 ;
        132:  q   <=  32'b00111100011000011011000010101010 ;
        133:  q   <=  32'b00111100011000110101111101110010 ;
        134:  q   <=  32'b00111100011001010000111000100001 ;
        135:  q   <=  32'b00111100011001101011110010110101 ;
        136:  q   <=  32'b00111100011010000110101100101111 ;
        137:  q   <=  32'b00111100011010100001100110001111 ;
        138:  q   <=  32'b00111100011010111100011111010101 ;
        139:  q   <=  32'b00111100011011010111011000000001 ;
        140:  q   <=  32'b00111100011011110010010000010011 ;
        141:  q   <=  32'b00111100011100001101001000001011 ;
        142:  q   <=  32'b00111100011100100111111111101001 ;
        143:  q   <=  32'b00111100011101000010110110101101 ;
        144:  q   <=  32'b00111100011101011101101101010111 ;
        145:  q   <=  32'b00111100011101111000100011100111 ;
        146:  q   <=  32'b00111100011110010011011001011110 ;
        147:  q   <=  32'b00111100011110101110001110111010 ;
        148:  q   <=  32'b00111100011111001001000011111100 ;
        149:  q   <=  32'b00111100011111100011111000100101 ;
        150:  q   <=  32'b00111100011111111110101100110100 ;
        151:  q   <=  32'b00111100100000001100110000010100 ;
        152:  q   <=  32'b00111100100000011010001010000010 ;
        153:  q   <=  32'b00111100100000100111100011100010 ;
        154:  q   <=  32'b00111100100000110100111100110110 ;
        155:  q   <=  32'b00111100100001000010010101111100 ;
        156:  q   <=  32'b00111100100001001111101110110110 ;
        157:  q   <=  32'b00111100100001011101000111100011 ;
        158:  q   <=  32'b00111100100001101010100000000011 ;
        159:  q   <=  32'b00111100100001110111111000010110 ;
        160:  q   <=  32'b00111100100010000101010000011101 ;
        161:  q   <=  32'b00111100100010010010101000010110 ;
        162:  q   <=  32'b00111100100010100000000000000011 ;
        163:  q   <=  32'b00111100100010101101010111100010 ;
        164:  q   <=  32'b00111100100010111010101110110101 ;
        165:  q   <=  32'b00111100100011001000000101111011 ;
        166:  q   <=  32'b00111100100011010101011100110100 ;
        167:  q   <=  32'b00111100100011100010110011100001 ;
        168:  q   <=  32'b00111100100011110000001010000000 ;
        169:  q   <=  32'b00111100100011111101100000010011 ;
        170:  q   <=  32'b00111100100100001010110110011001 ;
        171:  q   <=  32'b00111100100100011000001100010010 ;
        172:  q   <=  32'b00111100100100100101100001111110 ;
        173:  q   <=  32'b00111100100100110010110111011101 ;
        174:  q   <=  32'b00111100100101000000001100110000 ;
        175:  q   <=  32'b00111100100101001101100001110110 ;
        176:  q   <=  32'b00111100100101011010110110101111 ;
        177:  q   <=  32'b00111100100101101000001011011011 ;
        178:  q   <=  32'b00111100100101110101011111111011 ;
        179:  q   <=  32'b00111100100110000010110100001101 ;
        180:  q   <=  32'b00111100100110010000001000010011 ;
        181:  q   <=  32'b00111100100110011101011100001101 ;
        182:  q   <=  32'b00111100100110101010101111111001 ;
        183:  q   <=  32'b00111100100110111000000011011001 ;
        184:  q   <=  32'b00111100100111000101010110101100 ;
        185:  q   <=  32'b00111100100111010010101001110010 ;
        186:  q   <=  32'b00111100100111011111111100101100 ;
        187:  q   <=  32'b00111100100111101101001111011001 ;
        188:  q   <=  32'b00111100100111111010100001111001 ;
        189:  q   <=  32'b00111100101000000111110100001100 ;
        190:  q   <=  32'b00111100101000010101000110010011 ;
        191:  q   <=  32'b00111100101000100010011000001101 ;
        192:  q   <=  32'b00111100101000101111101001111010 ;
        193:  q   <=  32'b00111100101000111100111011011011 ;
        194:  q   <=  32'b00111100101001001010001100101111 ;
        195:  q   <=  32'b00111100101001010111011101110110 ;
        196:  q   <=  32'b00111100101001100100101110110001 ;
        197:  q   <=  32'b00111100101001110001111111011111 ;
        198:  q   <=  32'b00111100101001111111010000000000 ;
        199:  q   <=  32'b00111100101010001100100000010101 ;
        200:  q   <=  32'b00111100101010011001110000011101 ;
        201:  q   <=  32'b00111100101010100111000000011001 ;
        202:  q   <=  32'b00111100101010110100010000000111 ;
        203:  q   <=  32'b00111100101011000001011111101010 ;
        204:  q   <=  32'b00111100101011001110101110111111 ;
        205:  q   <=  32'b00111100101011011011111110001000 ;
        206:  q   <=  32'b00111100101011101001001101000101 ;
        207:  q   <=  32'b00111100101011110110011011110100 ;
        208:  q   <=  32'b00111100101100000011101010011000 ;
        209:  q   <=  32'b00111100101100010000111000101110 ;
        210:  q   <=  32'b00111100101100011110000110111000 ;
        211:  q   <=  32'b00111100101100101011010100110110 ;
        212:  q   <=  32'b00111100101100111000100010100110 ;
        213:  q   <=  32'b00111100101101000101110000001011 ;
        214:  q   <=  32'b00111100101101010010111101100010 ;
        215:  q   <=  32'b00111100101101100000001010101110 ;
        216:  q   <=  32'b00111100101101101101010111101100 ;
        217:  q   <=  32'b00111100101101111010100100011110 ;
        218:  q   <=  32'b00111100101110000111110001000100 ;
        219:  q   <=  32'b00111100101110010100111101011101 ;
        220:  q   <=  32'b00111100101110100010001001101010 ;
        221:  q   <=  32'b00111100101110101111010101101010 ;
        222:  q   <=  32'b00111100101110111100100001011101 ;
        223:  q   <=  32'b00111100101111001001101101000100 ;
        224:  q   <=  32'b00111100101111010110111000011110 ;
        225:  q   <=  32'b00111100101111100100000011101100 ;
        226:  q   <=  32'b00111100101111110001001110101110 ;
        227:  q   <=  32'b00111100101111111110011001100011 ;
        228:  q   <=  32'b00111100110000001011100100001100 ;
        229:  q   <=  32'b00111100110000011000101110101000 ;
        230:  q   <=  32'b00111100110000100101111000110111 ;
        231:  q   <=  32'b00111100110000110011000010111010 ;
        232:  q   <=  32'b00111100110001000000001100110001 ;
        233:  q   <=  32'b00111100110001001101010110011011 ;
        234:  q   <=  32'b00111100110001011010011111111001 ;
        235:  q   <=  32'b00111100110001100111101001001011 ;
        236:  q   <=  32'b00111100110001110100110010001111 ;
        237:  q   <=  32'b00111100110010000001111011001000 ;
        238:  q   <=  32'b00111100110010001111000011110100 ;
        239:  q   <=  32'b00111100110010011100001100010100 ;
        240:  q   <=  32'b00111100110010101001010100100111 ;
        241:  q   <=  32'b00111100110010110110011100101110 ;
        242:  q   <=  32'b00111100110011000011100100101000 ;
        243:  q   <=  32'b00111100110011010000101100010111 ;
        244:  q   <=  32'b00111100110011011101110011111000 ;
        245:  q   <=  32'b00111100110011101010111011001110 ;
        246:  q   <=  32'b00111100110011111000000010010111 ;
        247:  q   <=  32'b00111100110100000101001001010011 ;
        248:  q   <=  32'b00111100110100010010010000000011 ;
        249:  q   <=  32'b00111100110100011111010110100111 ;
        250:  q   <=  32'b00111100110100101100011100111111 ;
        251:  q   <=  32'b00111100110100111001100011001010 ;
        252:  q   <=  32'b00111100110101000110101001001001 ;
        253:  q   <=  32'b00111100110101010011101110111011 ;
        254:  q   <=  32'b00111100110101100000110100100001 ;
        255:  q   <=  32'b00111100110101101101111001111011 ;
        256:  q   <=  32'b00111100110101111010111111001001 ;
        257:  q   <=  32'b00111100110110001000000100001010 ;
        258:  q   <=  32'b00111100110110010101001000111111 ;
        259:  q   <=  32'b00111100110110100010001101101000 ;
        260:  q   <=  32'b00111100110110101111010010000100 ;
        261:  q   <=  32'b00111100110110111100010110010100 ;
        262:  q   <=  32'b00111100110111001001011010011000 ;
        263:  q   <=  32'b00111100110111010110011110001111 ;
        264:  q   <=  32'b00111100110111100011100001111010 ;
        265:  q   <=  32'b00111100110111110000100101011001 ;
        266:  q   <=  32'b00111100110111111101101000101100 ;
        267:  q   <=  32'b00111100111000001010101011110011 ;
        268:  q   <=  32'b00111100111000010111101110101101 ;
        269:  q   <=  32'b00111100111000100100110001011011 ;
        270:  q   <=  32'b00111100111000110001110011111100 ;
        271:  q   <=  32'b00111100111000111110110110010010 ;
        272:  q   <=  32'b00111100111001001011111000011011 ;
        273:  q   <=  32'b00111100111001011000111010011000 ;
        274:  q   <=  32'b00111100111001100101111100001001 ;
        275:  q   <=  32'b00111100111001110010111101101110 ;
        276:  q   <=  32'b00111100111001111111111111000110 ;
        277:  q   <=  32'b00111100111010001101000000010010 ;
        278:  q   <=  32'b00111100111010011010000001010010 ;
        279:  q   <=  32'b00111100111010100111000010000110 ;
        280:  q   <=  32'b00111100111010110100000010101110 ;
        281:  q   <=  32'b00111100111011000001000011001001 ;
        282:  q   <=  32'b00111100111011001110000011011000 ;
        283:  q   <=  32'b00111100111011011011000011011100 ;
        284:  q   <=  32'b00111100111011101000000011010010 ;
        285:  q   <=  32'b00111100111011110101000010111101 ;
        286:  q   <=  32'b00111100111100000010000010011100 ;
        287:  q   <=  32'b00111100111100001111000001101111 ;
        288:  q   <=  32'b00111100111100011100000000110101 ;
        289:  q   <=  32'b00111100111100101000111111101111 ;
        290:  q   <=  32'b00111100111100110101111110011101 ;
        291:  q   <=  32'b00111100111101000010111100111111 ;
        292:  q   <=  32'b00111100111101001111111011010101 ;
        293:  q   <=  32'b00111100111101011100111001011111 ;
        294:  q   <=  32'b00111100111101101001110111011101 ;
        295:  q   <=  32'b00111100111101110110110101001110 ;
        296:  q   <=  32'b00111100111110000011110010110100 ;
        297:  q   <=  32'b00111100111110010000110000001101 ;
        298:  q   <=  32'b00111100111110011101101101011010 ;
        299:  q   <=  32'b00111100111110101010101010011100 ;
        300:  q   <=  32'b00111100111110110111100111010001 ;
        301:  q   <=  32'b00111100111111000100100011111010 ;
        302:  q   <=  32'b00111100111111010001100000010111 ;
        303:  q   <=  32'b00111100111111011110011100101000 ;
        304:  q   <=  32'b00111100111111101011011000101101 ;
        305:  q   <=  32'b00111100111111111000010100100110 ;
        306:  q   <=  32'b00111101000000000010101000001001 ;
        307:  q   <=  32'b00111101000000001001000101111010 ;
        308:  q   <=  32'b00111101000000001111100011100100 ;
        309:  q   <=  32'b00111101000000010110000001001000 ;
        310:  q   <=  32'b00111101000000011100011110100111 ;
        311:  q   <=  32'b00111101000000100010111011111111 ;
        312:  q   <=  32'b00111101000000101001011001010010 ;
        313:  q   <=  32'b00111101000000101111110110011110 ;
        314:  q   <=  32'b00111101000000110110010011100100 ;
        315:  q   <=  32'b00111101000000111100110000100101 ;
        316:  q   <=  32'b00111101000001000011001101011111 ;
        317:  q   <=  32'b00111101000001001001101010010011 ;
        318:  q   <=  32'b00111101000001010000000111000010 ;
        319:  q   <=  32'b00111101000001010110100011101010 ;
        320:  q   <=  32'b00111101000001011101000000001101 ;
        321:  q   <=  32'b00111101000001100011011100101001 ;
        322:  q   <=  32'b00111101000001101001111001000000 ;
        323:  q   <=  32'b00111101000001110000010101010000 ;
        324:  q   <=  32'b00111101000001110110110001011011 ;
        325:  q   <=  32'b00111101000001111101001101011111 ;
        326:  q   <=  32'b00111101000010000011101001011110 ;
        327:  q   <=  32'b00111101000010001010000101010111 ;
        328:  q   <=  32'b00111101000010010000100001001001 ;
        329:  q   <=  32'b00111101000010010110111100110110 ;
        330:  q   <=  32'b00111101000010011101011000011101 ;
        331:  q   <=  32'b00111101000010100011110011111110 ;
        332:  q   <=  32'b00111101000010101010001111011001 ;
        333:  q   <=  32'b00111101000010110000101010101110 ;
        334:  q   <=  32'b00111101000010110111000101111101 ;
        335:  q   <=  32'b00111101000010111101100001000110 ;
        336:  q   <=  32'b00111101000011000011111100001001 ;
        337:  q   <=  32'b00111101000011001010010111000110 ;
        338:  q   <=  32'b00111101000011010000110001111101 ;
        339:  q   <=  32'b00111101000011010111001100101111 ;
        340:  q   <=  32'b00111101000011011101100111011010 ;
        341:  q   <=  32'b00111101000011100100000010000000 ;
        342:  q   <=  32'b00111101000011101010011100011111 ;
        343:  q   <=  32'b00111101000011110000110110111001 ;
        344:  q   <=  32'b00111101000011110111010001001100 ;
        345:  q   <=  32'b00111101000011111101101011011010 ;
        346:  q   <=  32'b00111101000100000100000101100010 ;
        347:  q   <=  32'b00111101000100001010011111100100 ;
        348:  q   <=  32'b00111101000100010000111001100000 ;
        349:  q   <=  32'b00111101000100010111010011010110 ;
        350:  q   <=  32'b00111101000100011101101101000111 ;
        351:  q   <=  32'b00111101000100100100000110110001 ;
        352:  q   <=  32'b00111101000100101010100000010110 ;
        353:  q   <=  32'b00111101000100110000111001110100 ;
        354:  q   <=  32'b00111101000100110111010011001101 ;
        355:  q   <=  32'b00111101000100111101101100100000 ;
        356:  q   <=  32'b00111101000101000100000101101101 ;
        357:  q   <=  32'b00111101000101001010011110110100 ;
        358:  q   <=  32'b00111101000101010000110111110101 ;
        359:  q   <=  32'b00111101000101010111010000110000 ;
        360:  q   <=  32'b00111101000101011101101001100110 ;
        361:  q   <=  32'b00111101000101100100000010010101 ;
        362:  q   <=  32'b00111101000101101010011010111111 ;
        363:  q   <=  32'b00111101000101110000110011100011 ;
        364:  q   <=  32'b00111101000101110111001100000001 ;
        365:  q   <=  32'b00111101000101111101100100011001 ;
        366:  q   <=  32'b00111101000110000011111100101011 ;
        367:  q   <=  32'b00111101000110001010010100110111 ;
        368:  q   <=  32'b00111101000110010000101100111110 ;
        369:  q   <=  32'b00111101000110010111000100111110 ;
        370:  q   <=  32'b00111101000110011101011100111001 ;
        371:  q   <=  32'b00111101000110100011110100101110 ;
        372:  q   <=  32'b00111101000110101010001100011101 ;
        373:  q   <=  32'b00111101000110110000100100000111 ;
        374:  q   <=  32'b00111101000110110110111011101010 ;
        375:  q   <=  32'b00111101000110111101010011001000 ;
        376:  q   <=  32'b00111101000111000011101010100000 ;
        377:  q   <=  32'b00111101000111001010000001110010 ;
        378:  q   <=  32'b00111101000111010000011000111110 ;
        379:  q   <=  32'b00111101000111010110110000000100 ;
        380:  q   <=  32'b00111101000111011101000111000100 ;
        381:  q   <=  32'b00111101000111100011011101111111 ;
        382:  q   <=  32'b00111101000111101001110100110100 ;
        383:  q   <=  32'b00111101000111110000001011100011 ;
        384:  q   <=  32'b00111101000111110110100010001100 ;
        385:  q   <=  32'b00111101000111111100111000110000 ;
        386:  q   <=  32'b00111101001000000011001111001101 ;
        387:  q   <=  32'b00111101001000001001100101100101 ;
        388:  q   <=  32'b00111101001000001111111011110111 ;
        389:  q   <=  32'b00111101001000010110010010000011 ;
        390:  q   <=  32'b00111101001000011100101000001010 ;
        391:  q   <=  32'b00111101001000100010111110001010 ;
        392:  q   <=  32'b00111101001000101001010100000101 ;
        393:  q   <=  32'b00111101001000101111101001111010 ;
        394:  q   <=  32'b00111101001000110101111111101010 ;
        395:  q   <=  32'b00111101001000111100010101010011 ;
        396:  q   <=  32'b00111101001001000010101010110111 ;
        397:  q   <=  32'b00111101001001001001000000010101 ;
        398:  q   <=  32'b00111101001001001111010101101101 ;
        399:  q   <=  32'b00111101001001010101101010111111 ;
        400:  q   <=  32'b00111101001001011100000000001100 ;
        401:  q   <=  32'b00111101001001100010010101010011 ;
        402:  q   <=  32'b00111101001001101000101010010100 ;
        403:  q   <=  32'b00111101001001101110111111001111 ;
        404:  q   <=  32'b00111101001001110101010100000101 ;
        405:  q   <=  32'b00111101001001111011101000110100 ;
        406:  q   <=  32'b00111101001010000001111101011110 ;
        407:  q   <=  32'b00111101001010001000010010000011 ;
        408:  q   <=  32'b00111101001010001110100110100001 ;
        409:  q   <=  32'b00111101001010010100111010111010 ;
        410:  q   <=  32'b00111101001010011011001111001101 ;
        411:  q   <=  32'b00111101001010100001100011011010 ;
        412:  q   <=  32'b00111101001010100111110111100010 ;
        413:  q   <=  32'b00111101001010101110001011100100 ;
        414:  q   <=  32'b00111101001010110100011111100000 ;
        415:  q   <=  32'b00111101001010111010110011010110 ;
        416:  q   <=  32'b00111101001011000001000111000111 ;
        417:  q   <=  32'b00111101001011000111011010110010 ;
        418:  q   <=  32'b00111101001011001101101110010111 ;
        419:  q   <=  32'b00111101001011010100000001110111 ;
        420:  q   <=  32'b00111101001011011010010101010000 ;
        421:  q   <=  32'b00111101001011100000101000100100 ;
        422:  q   <=  32'b00111101001011100110111011110011 ;
        423:  q   <=  32'b00111101001011101101001110111011 ;
        424:  q   <=  32'b00111101001011110011100001111110 ;
        425:  q   <=  32'b00111101001011111001110100111011 ;
        426:  q   <=  32'b00111101001100000000000111110011 ;
        427:  q   <=  32'b00111101001100000110011010100101 ;
        428:  q   <=  32'b00111101001100001100101101010001 ;
        429:  q   <=  32'b00111101001100010010111111110111 ;
        430:  q   <=  32'b00111101001100011001010010011000 ;
        431:  q   <=  32'b00111101001100011111100100110011 ;
        432:  q   <=  32'b00111101001100100101110111001000 ;
        433:  q   <=  32'b00111101001100101100001001011000 ;
        434:  q   <=  32'b00111101001100110010011011100010 ;
        435:  q   <=  32'b00111101001100111000101101100110 ;
        436:  q   <=  32'b00111101001100111110111111100101 ;
        437:  q   <=  32'b00111101001101000101010001011101 ;
        438:  q   <=  32'b00111101001101001011100011010001 ;
        439:  q   <=  32'b00111101001101010001110100111110 ;
        440:  q   <=  32'b00111101001101011000000110100110 ;
        441:  q   <=  32'b00111101001101011110011000001000 ;
        442:  q   <=  32'b00111101001101100100101001100101 ;
        443:  q   <=  32'b00111101001101101010111010111100 ;
        444:  q   <=  32'b00111101001101110001001100001101 ;
        445:  q   <=  32'b00111101001101110111011101011001 ;
        446:  q   <=  32'b00111101001101111101101110011111 ;
        447:  q   <=  32'b00111101001110000011111111011111 ;
        448:  q   <=  32'b00111101001110001010010000011010 ;
        449:  q   <=  32'b00111101001110010000100001001111 ;
        450:  q   <=  32'b00111101001110010110110001111110 ;
        451:  q   <=  32'b00111101001110011101000010101000 ;
        452:  q   <=  32'b00111101001110100011010011001100 ;
        453:  q   <=  32'b00111101001110101001100011101010 ;
        454:  q   <=  32'b00111101001110101111110100000011 ;
        455:  q   <=  32'b00111101001110110110000100010110 ;
        456:  q   <=  32'b00111101001110111100010100100100 ;
        457:  q   <=  32'b00111101001111000010100100101100 ;
        458:  q   <=  32'b00111101001111001000110100101110 ;
        459:  q   <=  32'b00111101001111001111000100101011 ;
        460:  q   <=  32'b00111101001111010101010100100010 ;
        461:  q   <=  32'b00111101001111011011100100010011 ;
        462:  q   <=  32'b00111101001111100001110011111111 ;
        463:  q   <=  32'b00111101001111101000000011100101 ;
        464:  q   <=  32'b00111101001111101110010011000110 ;
        465:  q   <=  32'b00111101001111110100100010100001 ;
        466:  q   <=  32'b00111101001111111010110001110110 ;
        467:  q   <=  32'b00111101010000000001000001000110 ;
        468:  q   <=  32'b00111101010000000111010000010000 ;
        469:  q   <=  32'b00111101010000001101011111010101 ;
        470:  q   <=  32'b00111101010000010011101110010100 ;
        471:  q   <=  32'b00111101010000011001111101001101 ;
        472:  q   <=  32'b00111101010000100000001100000001 ;
        473:  q   <=  32'b00111101010000100110011010101111 ;
        474:  q   <=  32'b00111101010000101100101001011000 ;
        475:  q   <=  32'b00111101010000110010110111111011 ;
        476:  q   <=  32'b00111101010000111001000110011000 ;
        477:  q   <=  32'b00111101010000111111010100110000 ;
        478:  q   <=  32'b00111101010001000101100011000011 ;
        479:  q   <=  32'b00111101010001001011110001001111 ;
        480:  q   <=  32'b00111101010001010001111111010110 ;
        481:  q   <=  32'b00111101010001011000001101011000 ;
        482:  q   <=  32'b00111101010001011110011011010100 ;
        483:  q   <=  32'b00111101010001100100101001001011 ;
        484:  q   <=  32'b00111101010001101010110110111100 ;
        485:  q   <=  32'b00111101010001110001000100100111 ;
        486:  q   <=  32'b00111101010001110111010010001101 ;
        487:  q   <=  32'b00111101010001111101011111101101 ;
        488:  q   <=  32'b00111101010010000011101101001000 ;
        489:  q   <=  32'b00111101010010001001111010011101 ;
        490:  q   <=  32'b00111101010010010000000111101101 ;
        491:  q   <=  32'b00111101010010010110010100110111 ;
        492:  q   <=  32'b00111101010010011100100001111011 ;
        493:  q   <=  32'b00111101010010100010101110111010 ;
        494:  q   <=  32'b00111101010010101000111011110100 ;
        495:  q   <=  32'b00111101010010101111001000101000 ;
        496:  q   <=  32'b00111101010010110101010101010110 ;
        497:  q   <=  32'b00111101010010111011100001111111 ;
        498:  q   <=  32'b00111101010011000001101110100010 ;
        499:  q   <=  32'b00111101010011000111111011000000 ;
        500:  q   <=  32'b00111101010011001110000111011000 ;
        501:  q   <=  32'b00111101010011010100010011101011 ;
        502:  q   <=  32'b00111101010011011010011111111000 ;
        503:  q   <=  32'b00111101010011100000101100000000 ;
        504:  q   <=  32'b00111101010011100110111000000010 ;
        505:  q   <=  32'b00111101010011101101000011111111 ;
        506:  q   <=  32'b00111101010011110011001111110110 ;
        507:  q   <=  32'b00111101010011111001011011101000 ;
        508:  q   <=  32'b00111101010011111111100111010100 ;
        509:  q   <=  32'b00111101010100000101110010111011 ;
        510:  q   <=  32'b00111101010100001011111110011100 ;
        511:  q   <=  32'b00111101010100010010001001111000 ;
        512:  q   <=  32'b00111101010100011000010101001110 ;
        513:  q   <=  32'b00111101010100011110100000011111 ;
        514:  q   <=  32'b00111101010100100100101011101010 ;
        515:  q   <=  32'b00111101010100101010110110110000 ;
        516:  q   <=  32'b00111101010100110001000001110000 ;
        517:  q   <=  32'b00111101010100110111001100101011 ;
        518:  q   <=  32'b00111101010100111101010111100000 ;
        519:  q   <=  32'b00111101010101000011100010010000 ;
        520:  q   <=  32'b00111101010101001001101100111011 ;
        521:  q   <=  32'b00111101010101001111110111100000 ;
        522:  q   <=  32'b00111101010101010110000001111111 ;
        523:  q   <=  32'b00111101010101011100001100011001 ;
        524:  q   <=  32'b00111101010101100010010110101101 ;
        525:  q   <=  32'b00111101010101101000100000111100 ;
        526:  q   <=  32'b00111101010101101110101011000110 ;
        527:  q   <=  32'b00111101010101110100110101001010 ;
        528:  q   <=  32'b00111101010101111010111111001001 ;
        529:  q   <=  32'b00111101010110000001001001000010 ;
        530:  q   <=  32'b00111101010110000111010010110110 ;
        531:  q   <=  32'b00111101010110001101011100100100 ;
        532:  q   <=  32'b00111101010110010011100110001101 ;
        533:  q   <=  32'b00111101010110011001101111110000 ;
        534:  q   <=  32'b00111101010110011111111001001110 ;
        535:  q   <=  32'b00111101010110100110000010100111 ;
        536:  q   <=  32'b00111101010110101100001011111010 ;
        537:  q   <=  32'b00111101010110110010010101001000 ;
        538:  q   <=  32'b00111101010110111000011110010000 ;
        539:  q   <=  32'b00111101010110111110100111010011 ;
        540:  q   <=  32'b00111101010111000100110000010000 ;
        541:  q   <=  32'b00111101010111001010111001001000 ;
        542:  q   <=  32'b00111101010111010001000001111011 ;
        543:  q   <=  32'b00111101010111010111001010101000 ;
        544:  q   <=  32'b00111101010111011101010011010000 ;
        545:  q   <=  32'b00111101010111100011011011110010 ;
        546:  q   <=  32'b00111101010111101001100100001111 ;
        547:  q   <=  32'b00111101010111101111101100100110 ;
        548:  q   <=  32'b00111101010111110101110100111000 ;
        549:  q   <=  32'b00111101010111111011111101000101 ;
        550:  q   <=  32'b00111101011000000010000101001100 ;
        551:  q   <=  32'b00111101011000001000001101001110 ;
        552:  q   <=  32'b00111101011000001110010101001011 ;
        553:  q   <=  32'b00111101011000010100011101000010 ;
        554:  q   <=  32'b00111101011000011010100100110011 ;
        555:  q   <=  32'b00111101011000100000101100100000 ;
        556:  q   <=  32'b00111101011000100110110100000111 ;
        557:  q   <=  32'b00111101011000101100111011101000 ;
        558:  q   <=  32'b00111101011000110011000011000100 ;
        559:  q   <=  32'b00111101011000111001001010011011 ;
        560:  q   <=  32'b00111101011000111111010001101100 ;
        561:  q   <=  32'b00111101011001000101011000111000 ;
        562:  q   <=  32'b00111101011001001011011111111111 ;
        563:  q   <=  32'b00111101011001010001100111000000 ;
        564:  q   <=  32'b00111101011001010111101101111100 ;
        565:  q   <=  32'b00111101011001011101110100110010 ;
        566:  q   <=  32'b00111101011001100011111011100100 ;
        567:  q   <=  32'b00111101011001101010000010001111 ;
        568:  q   <=  32'b00111101011001110000001000110110 ;
        569:  q   <=  32'b00111101011001110110001111010111 ;
        570:  q   <=  32'b00111101011001111100010101110010 ;
        571:  q   <=  32'b00111101011010000010011100001001 ;
        572:  q   <=  32'b00111101011010001000100010011010 ;
        573:  q   <=  32'b00111101011010001110101000100101 ;
        574:  q   <=  32'b00111101011010010100101110101100 ;
        575:  q   <=  32'b00111101011010011010110100101101 ;
        576:  q   <=  32'b00111101011010100000111010101000 ;
        577:  q   <=  32'b00111101011010100111000000011110 ;
        578:  q   <=  32'b00111101011010101101000110001111 ;
        579:  q   <=  32'b00111101011010110011001011111011 ;
        580:  q   <=  32'b00111101011010111001010001100001 ;
        581:  q   <=  32'b00111101011010111111010111000010 ;
        582:  q   <=  32'b00111101011011000101011100011110 ;
        583:  q   <=  32'b00111101011011001011100001110100 ;
        584:  q   <=  32'b00111101011011010001100111000101 ;
        585:  q   <=  32'b00111101011011010111101100010000 ;
        586:  q   <=  32'b00111101011011011101110001010111 ;
        587:  q   <=  32'b00111101011011100011110110011000 ;
        588:  q   <=  32'b00111101011011101001111011010011 ;
        589:  q   <=  32'b00111101011011110000000000001010 ;
        590:  q   <=  32'b00111101011011110110000100111011 ;
        591:  q   <=  32'b00111101011011111100001001100110 ;
        592:  q   <=  32'b00111101011100000010001110001101 ;
        593:  q   <=  32'b00111101011100001000010010101110 ;
        594:  q   <=  32'b00111101011100001110010111001010 ;
        595:  q   <=  32'b00111101011100010100011011100000 ;
        596:  q   <=  32'b00111101011100011010011111110001 ;
        597:  q   <=  32'b00111101011100100000100011111101 ;
        598:  q   <=  32'b00111101011100100110101000000100 ;
        599:  q   <=  32'b00111101011100101100101100000101 ;
        600:  q   <=  32'b00111101011100110010110000000001 ;
        601:  q   <=  32'b00111101011100111000110011111000 ;
        602:  q   <=  32'b00111101011100111110110111101010 ;
        603:  q   <=  32'b00111101011101000100111011010110 ;
        604:  q   <=  32'b00111101011101001010111110111101 ;
        605:  q   <=  32'b00111101011101010001000010011110 ;
        606:  q   <=  32'b00111101011101010111000101111011 ;
        607:  q   <=  32'b00111101011101011101001001010010 ;
        608:  q   <=  32'b00111101011101100011001100100011 ;
        609:  q   <=  32'b00111101011101101001001111110000 ;
        610:  q   <=  32'b00111101011101101111010010110111 ;
        611:  q   <=  32'b00111101011101110101010101111001 ;
        612:  q   <=  32'b00111101011101111011011000110110 ;
        613:  q   <=  32'b00111101011110000001011011101110 ;
        614:  q   <=  32'b00111101011110000111011110100000 ;
        615:  q   <=  32'b00111101011110001101100001001101 ;
        616:  q   <=  32'b00111101011110010011100011110100 ;
        617:  q   <=  32'b00111101011110011001100110010111 ;
        618:  q   <=  32'b00111101011110011111101000110100 ;
        619:  q   <=  32'b00111101011110100101101011001100 ;
        620:  q   <=  32'b00111101011110101011101101011111 ;
        621:  q   <=  32'b00111101011110110001101111101100 ;
        622:  q   <=  32'b00111101011110110111110001110101 ;
        623:  q   <=  32'b00111101011110111101110011111000 ;
        624:  q   <=  32'b00111101011111000011110101110101 ;
        625:  q   <=  32'b00111101011111001001110111101110 ;
        626:  q   <=  32'b00111101011111001111111001100001 ;
        627:  q   <=  32'b00111101011111010101111011001111 ;
        628:  q   <=  32'b00111101011111011011111100111000 ;
        629:  q   <=  32'b00111101011111100001111110011100 ;
        630:  q   <=  32'b00111101011111100111111111111010 ;
        631:  q   <=  32'b00111101011111101110000001010011 ;
        632:  q   <=  32'b00111101011111110100000010100111 ;
        633:  q   <=  32'b00111101011111111010000011110110 ;
        634:  q   <=  32'b00111101100000000000000010100000 ;
        635:  q   <=  32'b00111101100000000011000011000010 ;
        636:  q   <=  32'b00111101100000000110000011100001 ;
        637:  q   <=  32'b00111101100000001001000011111110 ;
        638:  q   <=  32'b00111101100000001100000100011001 ;
        639:  q   <=  32'b00111101100000001111000100110000 ;
        640:  q   <=  32'b00111101100000010010000101000110 ;
        641:  q   <=  32'b00111101100000010101000101011000 ;
        642:  q   <=  32'b00111101100000011000000101101000 ;
        643:  q   <=  32'b00111101100000011011000101110101 ;
        644:  q   <=  32'b00111101100000011110000110000000 ;
        645:  q   <=  32'b00111101100000100001000110001000 ;
        646:  q   <=  32'b00111101100000100100000110001110 ;
        647:  q   <=  32'b00111101100000100111000110010001 ;
        648:  q   <=  32'b00111101100000101010000110010001 ;
        649:  q   <=  32'b00111101100000101101000110001111 ;
        650:  q   <=  32'b00111101100000110000000110001010 ;
        651:  q   <=  32'b00111101100000110011000110000011 ;
        652:  q   <=  32'b00111101100000110110000101111001 ;
        653:  q   <=  32'b00111101100000111001000101101101 ;
        654:  q   <=  32'b00111101100000111100000101011101 ;
        655:  q   <=  32'b00111101100000111111000101001100 ;
        656:  q   <=  32'b00111101100001000010000100110111 ;
        657:  q   <=  32'b00111101100001000101000100100001 ;
        658:  q   <=  32'b00111101100001001000000100000111 ;
        659:  q   <=  32'b00111101100001001011000011101011 ;
        660:  q   <=  32'b00111101100001001110000011001100 ;
        661:  q   <=  32'b00111101100001010001000010101011 ;
        662:  q   <=  32'b00111101100001010100000010000111 ;
        663:  q   <=  32'b00111101100001010111000001100001 ;
        664:  q   <=  32'b00111101100001011010000000111000 ;
        665:  q   <=  32'b00111101100001011101000000001101 ;
        666:  q   <=  32'b00111101100001011111111111011111 ;
        667:  q   <=  32'b00111101100001100010111110101110 ;
        668:  q   <=  32'b00111101100001100101111101111011 ;
        669:  q   <=  32'b00111101100001101000111101000101 ;
        670:  q   <=  32'b00111101100001101011111100001101 ;
        671:  q   <=  32'b00111101100001101110111011010010 ;
        672:  q   <=  32'b00111101100001110001111010010100 ;
        673:  q   <=  32'b00111101100001110100111001010100 ;
        674:  q   <=  32'b00111101100001110111111000010010 ;
        675:  q   <=  32'b00111101100001111010110111001101 ;
        676:  q   <=  32'b00111101100001111101110110000101 ;
        677:  q   <=  32'b00111101100010000000110100111011 ;
        678:  q   <=  32'b00111101100010000011110011101110 ;
        679:  q   <=  32'b00111101100010000110110010011110 ;
        680:  q   <=  32'b00111101100010001001110001001101 ;
        681:  q   <=  32'b00111101100010001100101111111000 ;
        682:  q   <=  32'b00111101100010001111101110100001 ;
        683:  q   <=  32'b00111101100010010010101101000111 ;
        684:  q   <=  32'b00111101100010010101101011101011 ;
        685:  q   <=  32'b00111101100010011000101010001100 ;
        686:  q   <=  32'b00111101100010011011101000101011 ;
        687:  q   <=  32'b00111101100010011110100111000111 ;
        688:  q   <=  32'b00111101100010100001100101100001 ;
        689:  q   <=  32'b00111101100010100100100011111000 ;
        690:  q   <=  32'b00111101100010100111100010001101 ;
        691:  q   <=  32'b00111101100010101010100000011111 ;
        692:  q   <=  32'b00111101100010101101011110101110 ;
        693:  q   <=  32'b00111101100010110000011100111011 ;
        694:  q   <=  32'b00111101100010110011011011000101 ;
        695:  q   <=  32'b00111101100010110110011001001101 ;
        696:  q   <=  32'b00111101100010111001010111010011 ;
        697:  q   <=  32'b00111101100010111100010101010101 ;
        698:  q   <=  32'b00111101100010111111010011010110 ;
        699:  q   <=  32'b00111101100011000010010001010011 ;
        700:  q   <=  32'b00111101100011000101001111001110 ;
        701:  q   <=  32'b00111101100011001000001101000111 ;
        702:  q   <=  32'b00111101100011001011001010111101 ;
        703:  q   <=  32'b00111101100011001110001000110001 ;
        704:  q   <=  32'b00111101100011010001000110100010 ;
        705:  q   <=  32'b00111101100011010100000100010000 ;
        706:  q   <=  32'b00111101100011010111000001111100 ;
        707:  q   <=  32'b00111101100011011001111111100110 ;
        708:  q   <=  32'b00111101100011011100111101001100 ;
        709:  q   <=  32'b00111101100011011111111010110001 ;
        710:  q   <=  32'b00111101100011100010111000010011 ;
        711:  q   <=  32'b00111101100011100101110101110010 ;
        712:  q   <=  32'b00111101100011101000110011001111 ;
        713:  q   <=  32'b00111101100011101011110000101001 ;
        714:  q   <=  32'b00111101100011101110101110000001 ;
        715:  q   <=  32'b00111101100011110001101011010110 ;
        716:  q   <=  32'b00111101100011110100101000101001 ;
        717:  q   <=  32'b00111101100011110111100101111001 ;
        718:  q   <=  32'b00111101100011111010100011000111 ;
        719:  q   <=  32'b00111101100011111101100000010010 ;
        720:  q   <=  32'b00111101100100000000011101011011 ;
        721:  q   <=  32'b00111101100100000011011010100001 ;
        722:  q   <=  32'b00111101100100000110010111100100 ;
        723:  q   <=  32'b00111101100100001001010100100110 ;
        724:  q   <=  32'b00111101100100001100010001100100 ;
        725:  q   <=  32'b00111101100100001111001110100000 ;
        726:  q   <=  32'b00111101100100010010001011011010 ;
        727:  q   <=  32'b00111101100100010101001000010001 ;
        728:  q   <=  32'b00111101100100011000000101000110 ;
        729:  q   <=  32'b00111101100100011011000001111000 ;
        730:  q   <=  32'b00111101100100011101111110100111 ;
        731:  q   <=  32'b00111101100100100000111011010100 ;
        732:  q   <=  32'b00111101100100100011110111111111 ;
        733:  q   <=  32'b00111101100100100110110100100111 ;
        734:  q   <=  32'b00111101100100101001110001001101 ;
        735:  q   <=  32'b00111101100100101100101101110000 ;
        736:  q   <=  32'b00111101100100101111101010010000 ;
        737:  q   <=  32'b00111101100100110010100110101110 ;
        738:  q   <=  32'b00111101100100110101100011001010 ;
        739:  q   <=  32'b00111101100100111000011111100011 ;
        740:  q   <=  32'b00111101100100111011011011111010 ;
        741:  q   <=  32'b00111101100100111110011000001110 ;
        742:  q   <=  32'b00111101100101000001010100011111 ;
        743:  q   <=  32'b00111101100101000100010000101110 ;
        744:  q   <=  32'b00111101100101000111001100111011 ;
        745:  q   <=  32'b00111101100101001010001001000101 ;
        746:  q   <=  32'b00111101100101001101000101001101 ;
        747:  q   <=  32'b00111101100101010000000001010010 ;
        748:  q   <=  32'b00111101100101010010111101010101 ;
        749:  q   <=  32'b00111101100101010101111001010101 ;
        750:  q   <=  32'b00111101100101011000110101010011 ;
        751:  q   <=  32'b00111101100101011011110001001110 ;
        752:  q   <=  32'b00111101100101011110101101000111 ;
        753:  q   <=  32'b00111101100101100001101000111101 ;
        754:  q   <=  32'b00111101100101100100100100110001 ;
        755:  q   <=  32'b00111101100101100111100000100010 ;
        756:  q   <=  32'b00111101100101101010011100010001 ;
        757:  q   <=  32'b00111101100101101101010111111101 ;
        758:  q   <=  32'b00111101100101110000010011100111 ;
        759:  q   <=  32'b00111101100101110011001111001111 ;
        760:  q   <=  32'b00111101100101110110001010110100 ;
        761:  q   <=  32'b00111101100101111001000110010110 ;
        762:  q   <=  32'b00111101100101111100000001110110 ;
        763:  q   <=  32'b00111101100101111110111101010100 ;
        764:  q   <=  32'b00111101100110000001111000101111 ;
        765:  q   <=  32'b00111101100110000100110100000111 ;
        766:  q   <=  32'b00111101100110000111101111011101 ;
        767:  q   <=  32'b00111101100110001010101010110001 ;
        768:  q   <=  32'b00111101100110001101100110000010 ;
        769:  q   <=  32'b00111101100110010000100001010001 ;
        770:  q   <=  32'b00111101100110010011011100011101 ;
        771:  q   <=  32'b00111101100110010110010111100111 ;
        772:  q   <=  32'b00111101100110011001010010101110 ;
        773:  q   <=  32'b00111101100110011100001101110011 ;
        774:  q   <=  32'b00111101100110011111001000110110 ;
        775:  q   <=  32'b00111101100110100010000011110110 ;
        776:  q   <=  32'b00111101100110100100111110110011 ;
        777:  q   <=  32'b00111101100110100111111001101110 ;
        778:  q   <=  32'b00111101100110101010110100100111 ;
        779:  q   <=  32'b00111101100110101101101111011101 ;
        780:  q   <=  32'b00111101100110110000101010010001 ;
        781:  q   <=  32'b00111101100110110011100101000010 ;
        782:  q   <=  32'b00111101100110110110011111110001 ;
        783:  q   <=  32'b00111101100110111001011010011101 ;
        784:  q   <=  32'b00111101100110111100010101000111 ;
        785:  q   <=  32'b00111101100110111111001111101110 ;
        786:  q   <=  32'b00111101100111000010001010010011 ;
        787:  q   <=  32'b00111101100111000101000100110110 ;
        788:  q   <=  32'b00111101100111000111111111010110 ;
        789:  q   <=  32'b00111101100111001010111001110100 ;
        790:  q   <=  32'b00111101100111001101110100001111 ;
        791:  q   <=  32'b00111101100111010000101110101000 ;
        792:  q   <=  32'b00111101100111010011101000111110 ;
        793:  q   <=  32'b00111101100111010110100011010010 ;
        794:  q   <=  32'b00111101100111011001011101100100 ;
        795:  q   <=  32'b00111101100111011100010111110011 ;
        796:  q   <=  32'b00111101100111011111010001111111 ;
        797:  q   <=  32'b00111101100111100010001100001001 ;
        798:  q   <=  32'b00111101100111100101000110010001 ;
        799:  q   <=  32'b00111101100111101000000000010110 ;
        800:  q   <=  32'b00111101100111101010111010011001 ;
        801:  q   <=  32'b00111101100111101101110100011010 ;
        802:  q   <=  32'b00111101100111110000101110011000 ;
        803:  q   <=  32'b00111101100111110011101000010011 ;
        804:  q   <=  32'b00111101100111110110100010001100 ;
        805:  q   <=  32'b00111101100111111001011100000011 ;
        806:  q   <=  32'b00111101100111111100010101110111 ;
        807:  q   <=  32'b00111101100111111111001111101001 ;
        808:  q   <=  32'b00111101101000000010001001011001 ;
        809:  q   <=  32'b00111101101000000101000011000110 ;
        810:  q   <=  32'b00111101101000000111111100110000 ;
        811:  q   <=  32'b00111101101000001010110110011000 ;
        812:  q   <=  32'b00111101101000001101101111111110 ;
        813:  q   <=  32'b00111101101000010000101001100001 ;
        814:  q   <=  32'b00111101101000010011100011000010 ;
        815:  q   <=  32'b00111101101000010110011100100001 ;
        816:  q   <=  32'b00111101101000011001010101111101 ;
        817:  q   <=  32'b00111101101000011100001111010111 ;
        818:  q   <=  32'b00111101101000011111001000101110 ;
        819:  q   <=  32'b00111101101000100010000010000011 ;
        820:  q   <=  32'b00111101101000100100111011010101 ;
        821:  q   <=  32'b00111101101000100111110100100101 ;
        822:  q   <=  32'b00111101101000101010101101110011 ;
        823:  q   <=  32'b00111101101000101101100110111110 ;
        824:  q   <=  32'b00111101101000110000100000000111 ;
        825:  q   <=  32'b00111101101000110011011001001101 ;
        826:  q   <=  32'b00111101101000110110010010010001 ;
        827:  q   <=  32'b00111101101000111001001011010010 ;
        828:  q   <=  32'b00111101101000111100000100010010 ;
        829:  q   <=  32'b00111101101000111110111101001110 ;
        830:  q   <=  32'b00111101101001000001110110001001 ;
        831:  q   <=  32'b00111101101001000100101111000001 ;
        832:  q   <=  32'b00111101101001000111100111110110 ;
        833:  q   <=  32'b00111101101001001010100000101001 ;
        834:  q   <=  32'b00111101101001001101011001011010 ;
        835:  q   <=  32'b00111101101001010000010010001000 ;
        836:  q   <=  32'b00111101101001010011001010110100 ;
        837:  q   <=  32'b00111101101001010110000011011110 ;
        838:  q   <=  32'b00111101101001011000111100000101 ;
        839:  q   <=  32'b00111101101001011011110100101010 ;
        840:  q   <=  32'b00111101101001011110101101001100 ;
        841:  q   <=  32'b00111101101001100001100101101100 ;
        842:  q   <=  32'b00111101101001100100011110001010 ;
        843:  q   <=  32'b00111101101001100111010110100101 ;
        844:  q   <=  32'b00111101101001101010001110111110 ;
        845:  q   <=  32'b00111101101001101101000111010100 ;
        846:  q   <=  32'b00111101101001101111111111101000 ;
        847:  q   <=  32'b00111101101001110010110111111010 ;
        848:  q   <=  32'b00111101101001110101110000001001 ;
        849:  q   <=  32'b00111101101001111000101000010110 ;
        850:  q   <=  32'b00111101101001111011100000100000 ;
        851:  q   <=  32'b00111101101001111110011000101000 ;
        852:  q   <=  32'b00111101101010000001010000101110 ;
        853:  q   <=  32'b00111101101010000100001000110001 ;
        854:  q   <=  32'b00111101101010000111000000110010 ;
        855:  q   <=  32'b00111101101010001001111000110001 ;
        856:  q   <=  32'b00111101101010001100110000101101 ;
        857:  q   <=  32'b00111101101010001111101000100111 ;
        858:  q   <=  32'b00111101101010010010100000011110 ;
        859:  q   <=  32'b00111101101010010101011000010011 ;
        860:  q   <=  32'b00111101101010011000010000000110 ;
        861:  q   <=  32'b00111101101010011011000111110110 ;
        862:  q   <=  32'b00111101101010011101111111100100 ;
        863:  q   <=  32'b00111101101010100000110111010000 ;
        864:  q   <=  32'b00111101101010100011101110111001 ;
        865:  q   <=  32'b00111101101010100110100110100000 ;
        866:  q   <=  32'b00111101101010101001011110000100 ;
        867:  q   <=  32'b00111101101010101100010101100110 ;
        868:  q   <=  32'b00111101101010101111001101000110 ;
        869:  q   <=  32'b00111101101010110010000100100100 ;
        870:  q   <=  32'b00111101101010110100111011111111 ;
        871:  q   <=  32'b00111101101010110111110011010111 ;
        872:  q   <=  32'b00111101101010111010101010101101 ;
        873:  q   <=  32'b00111101101010111101100010000001 ;
        874:  q   <=  32'b00111101101011000000011001010011 ;
        875:  q   <=  32'b00111101101011000011010000100010 ;
        876:  q   <=  32'b00111101101011000110000111101111 ;
        877:  q   <=  32'b00111101101011001000111110111001 ;
        878:  q   <=  32'b00111101101011001011110110000010 ;
        879:  q   <=  32'b00111101101011001110101101000111 ;
        880:  q   <=  32'b00111101101011010001100100001011 ;
        881:  q   <=  32'b00111101101011010100011011001100 ;
        882:  q   <=  32'b00111101101011010111010010001010 ;
        883:  q   <=  32'b00111101101011011010001001000111 ;
        884:  q   <=  32'b00111101101011011101000000000001 ;
        885:  q   <=  32'b00111101101011011111110110111000 ;
        886:  q   <=  32'b00111101101011100010101101101110 ;
        887:  q   <=  32'b00111101101011100101100100100001 ;
        888:  q   <=  32'b00111101101011101000011011010001 ;
        889:  q   <=  32'b00111101101011101011010010000000 ;
        890:  q   <=  32'b00111101101011101110001000101100 ;
        891:  q   <=  32'b00111101101011110000111111010101 ;
        892:  q   <=  32'b00111101101011110011110101111100 ;
        893:  q   <=  32'b00111101101011110110101100100001 ;
        894:  q   <=  32'b00111101101011111001100011000100 ;
        895:  q   <=  32'b00111101101011111100011001100100 ;
        896:  q   <=  32'b00111101101011111111010000000010 ;
        897:  q   <=  32'b00111101101100000010000110011101 ;
        898:  q   <=  32'b00111101101100000100111100110110 ;
        899:  q   <=  32'b00111101101100000111110011001101 ;
        900:  q   <=  32'b00111101101100001010101001100010 ;
        901:  q   <=  32'b00111101101100001101011111110100 ;
        902:  q   <=  32'b00111101101100010000010110000100 ;
        903:  q   <=  32'b00111101101100010011001100010001 ;
        904:  q   <=  32'b00111101101100010110000010011100 ;
        905:  q   <=  32'b00111101101100011000111000100101 ;
        906:  q   <=  32'b00111101101100011011101110101100 ;
        907:  q   <=  32'b00111101101100011110100100110000 ;
        908:  q   <=  32'b00111101101100100001011010110010 ;
        909:  q   <=  32'b00111101101100100100010000110001 ;
        910:  q   <=  32'b00111101101100100111000110101111 ;
        911:  q   <=  32'b00111101101100101001111100101001 ;
        912:  q   <=  32'b00111101101100101100110010100010 ;
        913:  q   <=  32'b00111101101100101111101000011000 ;
        914:  q   <=  32'b00111101101100110010011110001100 ;
        915:  q   <=  32'b00111101101100110101010011111110 ;
        916:  q   <=  32'b00111101101100111000001001101101 ;
        917:  q   <=  32'b00111101101100111010111111011010 ;
        918:  q   <=  32'b00111101101100111101110101000100 ;
        919:  q   <=  32'b00111101101101000000101010101101 ;
        920:  q   <=  32'b00111101101101000011100000010011 ;
        921:  q   <=  32'b00111101101101000110010101110110 ;
        922:  q   <=  32'b00111101101101001001001011011000 ;
        923:  q   <=  32'b00111101101101001100000000110111 ;
        924:  q   <=  32'b00111101101101001110110110010011 ;
        925:  q   <=  32'b00111101101101010001101011101110 ;
        926:  q   <=  32'b00111101101101010100100001000110 ;
        927:  q   <=  32'b00111101101101010111010110011100 ;
        928:  q   <=  32'b00111101101101011010001011101111 ;
        929:  q   <=  32'b00111101101101011101000001000000 ;
        930:  q   <=  32'b00111101101101011111110110001111 ;
        931:  q   <=  32'b00111101101101100010101011011100 ;
        932:  q   <=  32'b00111101101101100101100000100110 ;
        933:  q   <=  32'b00111101101101101000010101101110 ;
        934:  q   <=  32'b00111101101101101011001010110100 ;
        935:  q   <=  32'b00111101101101101101111111110111 ;
        936:  q   <=  32'b00111101101101110000110100111000 ;
        937:  q   <=  32'b00111101101101110011101001110111 ;
        938:  q   <=  32'b00111101101101110110011110110011 ;
        939:  q   <=  32'b00111101101101111001010011101101 ;
        940:  q   <=  32'b00111101101101111100001000100101 ;
        941:  q   <=  32'b00111101101101111110111101011010 ;
        942:  q   <=  32'b00111101101110000001110010001110 ;
        943:  q   <=  32'b00111101101110000100100110111111 ;
        944:  q   <=  32'b00111101101110000111011011101101 ;
        945:  q   <=  32'b00111101101110001010010000011010 ;
        946:  q   <=  32'b00111101101110001101000101000100 ;
        947:  q   <=  32'b00111101101110001111111001101011 ;
        948:  q   <=  32'b00111101101110010010101110010001 ;
        949:  q   <=  32'b00111101101110010101100010110100 ;
        950:  q   <=  32'b00111101101110011000010111010101 ;
        951:  q   <=  32'b00111101101110011011001011110011 ;
        952:  q   <=  32'b00111101101110011110000000010000 ;
        953:  q   <=  32'b00111101101110100000110100101010 ;
        954:  q   <=  32'b00111101101110100011101001000001 ;
        955:  q   <=  32'b00111101101110100110011101010111 ;
        956:  q   <=  32'b00111101101110101001010001101010 ;
        957:  q   <=  32'b00111101101110101100000101111011 ;
        958:  q   <=  32'b00111101101110101110111010001001 ;
        959:  q   <=  32'b00111101101110110001101110010110 ;
        960:  q   <=  32'b00111101101110110100100010100000 ;
        961:  q   <=  32'b00111101101110110111010110101000 ;
        962:  q   <=  32'b00111101101110111010001010101101 ;
        963:  q   <=  32'b00111101101110111100111110110000 ;
        964:  q   <=  32'b00111101101110111111110010110001 ;
        965:  q   <=  32'b00111101101111000010100110110000 ;
        966:  q   <=  32'b00111101101111000101011010101100 ;
        967:  q   <=  32'b00111101101111001000001110100110 ;
        968:  q   <=  32'b00111101101111001011000010011110 ;
        969:  q   <=  32'b00111101101111001101110110010011 ;
        970:  q   <=  32'b00111101101111010000101010000111 ;
        971:  q   <=  32'b00111101101111010011011101111000 ;
        972:  q   <=  32'b00111101101111010110010001100110 ;
        973:  q   <=  32'b00111101101111011001000101010011 ;
        974:  q   <=  32'b00111101101111011011111000111101 ;
        975:  q   <=  32'b00111101101111011110101100100101 ;
        976:  q   <=  32'b00111101101111100001100000001011 ;
        977:  q   <=  32'b00111101101111100100010011101110 ;
        978:  q   <=  32'b00111101101111100111000111001111 ;
        979:  q   <=  32'b00111101101111101001111010101110 ;
        980:  q   <=  32'b00111101101111101100101110001011 ;
        981:  q   <=  32'b00111101101111101111100001100101 ;
        982:  q   <=  32'b00111101101111110010010100111101 ;
        983:  q   <=  32'b00111101101111110101001000010011 ;
        984:  q   <=  32'b00111101101111110111111011100110 ;
        985:  q   <=  32'b00111101101111111010101110111000 ;
        986:  q   <=  32'b00111101101111111101100010000111 ;
        987:  q   <=  32'b00111101110000000000010101010011 ;
        988:  q   <=  32'b00111101110000000011001000011110 ;
        989:  q   <=  32'b00111101110000000101111011100110 ;
        990:  q   <=  32'b00111101110000001000101110101100 ;
        991:  q   <=  32'b00111101110000001011100001110000 ;
        992:  q   <=  32'b00111101110000001110010100110001 ;
        993:  q   <=  32'b00111101110000010001000111110001 ;
        994:  q   <=  32'b00111101110000010011111010101110 ;
        995:  q   <=  32'b00111101110000010110101101101000 ;
        996:  q   <=  32'b00111101110000011001100000100001 ;
        997:  q   <=  32'b00111101110000011100010011010111 ;
        998:  q   <=  32'b00111101110000011111000110001011 ;
        999:  q   <=  32'b00111101110000100001111000111101 ;
        1000:  q   <=  32'b00111101110000100100101011101100 ;
        1001:  q   <=  32'b00111101110000100111011110011010 ;
        1002:  q   <=  32'b00111101110000101010010001000101 ;
        1003:  q   <=  32'b00111101110000101101000011101101 ;
        1004:  q   <=  32'b00111101110000101111110110010100 ;
        1005:  q   <=  32'b00111101110000110010101000111000 ;
        1006:  q   <=  32'b00111101110000110101011011011010 ;
        1007:  q   <=  32'b00111101110000111000001101111010 ;
        1008:  q   <=  32'b00111101110000111011000000011000 ;
        1009:  q   <=  32'b00111101110000111101110010110011 ;
        1010:  q   <=  32'b00111101110001000000100101001100 ;
        1011:  q   <=  32'b00111101110001000011010111100011 ;
        1012:  q   <=  32'b00111101110001000110001001111000 ;
        1013:  q   <=  32'b00111101110001001000111100001010 ;
        1014:  q   <=  32'b00111101110001001011101110011010 ;
        1015:  q   <=  32'b00111101110001001110100000101000 ;
        1016:  q   <=  32'b00111101110001010001010010110100 ;
        1017:  q   <=  32'b00111101110001010100000100111101 ;
        1018:  q   <=  32'b00111101110001010110110111000101 ;
        1019:  q   <=  32'b00111101110001011001101001001010 ;
        1020:  q   <=  32'b00111101110001011100011011001100 ;
        1021:  q   <=  32'b00111101110001011111001101001101 ;
        1022:  q   <=  32'b00111101110001100001111111001011 ;
        1023:  q   <=  32'b00111101110001100100110001000111 ;
        1024:  q   <=  32'b00111101110001100111100011000001 ;
        1025:  q   <=  32'b00111101110001101010010100111001 ;
        1026:  q   <=  32'b00111101110001101101000110101110 ;
        1027:  q   <=  32'b00111101110001101111111000100010 ;
        1028:  q   <=  32'b00111101110001110010101010010011 ;
        1029:  q   <=  32'b00111101110001110101011100000001 ;
        1030:  q   <=  32'b00111101110001111000001101101110 ;
        1031:  q   <=  32'b00111101110001111010111111011000 ;
        1032:  q   <=  32'b00111101110001111101110001000000 ;
        1033:  q   <=  32'b00111101110010000000100010100110 ;
        1034:  q   <=  32'b00111101110010000011010100001010 ;
        1035:  q   <=  32'b00111101110010000110000101101011 ;
        1036:  q   <=  32'b00111101110010001000110111001011 ;
        1037:  q   <=  32'b00111101110010001011101000101000 ;
        1038:  q   <=  32'b00111101110010001110011010000011 ;
        1039:  q   <=  32'b00111101110010010001001011011011 ;
        1040:  q   <=  32'b00111101110010010011111100110010 ;
        1041:  q   <=  32'b00111101110010010110101110000110 ;
        1042:  q   <=  32'b00111101110010011001011111011000 ;
        1043:  q   <=  32'b00111101110010011100010000101000 ;
        1044:  q   <=  32'b00111101110010011111000001110101 ;
        1045:  q   <=  32'b00111101110010100001110011000000 ;
        1046:  q   <=  32'b00111101110010100100100100001010 ;
        1047:  q   <=  32'b00111101110010100111010101010001 ;
        1048:  q   <=  32'b00111101110010101010000110010101 ;
        1049:  q   <=  32'b00111101110010101100110111011000 ;
        1050:  q   <=  32'b00111101110010101111101000011000 ;
        1051:  q   <=  32'b00111101110010110010011001010110 ;
        1052:  q   <=  32'b00111101110010110101001010010010 ;
        1053:  q   <=  32'b00111101110010110111111011001100 ;
        1054:  q   <=  32'b00111101110010111010101100000100 ;
        1055:  q   <=  32'b00111101110010111101011100111001 ;
        1056:  q   <=  32'b00111101110011000000001101101100 ;
        1057:  q   <=  32'b00111101110011000010111110011101 ;
        1058:  q   <=  32'b00111101110011000101101111001100 ;
        1059:  q   <=  32'b00111101110011001000011111111000 ;
        1060:  q   <=  32'b00111101110011001011010000100011 ;
        1061:  q   <=  32'b00111101110011001110000001001011 ;
        1062:  q   <=  32'b00111101110011010000110001110001 ;
        1063:  q   <=  32'b00111101110011010011100010010101 ;
        1064:  q   <=  32'b00111101110011010110010010110110 ;
        1065:  q   <=  32'b00111101110011011001000011010110 ;
        1066:  q   <=  32'b00111101110011011011110011110011 ;
        1067:  q   <=  32'b00111101110011011110100100001110 ;
        1068:  q   <=  32'b00111101110011100001010100100111 ;
        1069:  q   <=  32'b00111101110011100100000100111110 ;
        1070:  q   <=  32'b00111101110011100110110101010010 ;
        1071:  q   <=  32'b00111101110011101001100101100100 ;
        1072:  q   <=  32'b00111101110011101100010101110101 ;
        1073:  q   <=  32'b00111101110011101111000110000010 ;
        1074:  q   <=  32'b00111101110011110001110110001110 ;
        1075:  q   <=  32'b00111101110011110100100110011000 ;
        1076:  q   <=  32'b00111101110011110111010110011111 ;
        1077:  q   <=  32'b00111101110011111010000110100100 ;
        1078:  q   <=  32'b00111101110011111100110110100111 ;
        1079:  q   <=  32'b00111101110011111111100110101000 ;
        1080:  q   <=  32'b00111101110100000010010110100111 ;
        1081:  q   <=  32'b00111101110100000101000110100011 ;
        1082:  q   <=  32'b00111101110100000111110110011110 ;
        1083:  q   <=  32'b00111101110100001010100110010110 ;
        1084:  q   <=  32'b00111101110100001101010110001100 ;
        1085:  q   <=  32'b00111101110100010000000110000000 ;
        1086:  q   <=  32'b00111101110100010010110101110001 ;
        1087:  q   <=  32'b00111101110100010101100101100001 ;
        1088:  q   <=  32'b00111101110100011000010101001110 ;
        1089:  q   <=  32'b00111101110100011011000100111001 ;
        1090:  q   <=  32'b00111101110100011101110100100010 ;
        1091:  q   <=  32'b00111101110100100000100100001001 ;
        1092:  q   <=  32'b00111101110100100011010011101110 ;
        1093:  q   <=  32'b00111101110100100110000011010000 ;
        1094:  q   <=  32'b00111101110100101000110010110000 ;
        1095:  q   <=  32'b00111101110100101011100010001111 ;
        1096:  q   <=  32'b00111101110100101110010001101011 ;
        1097:  q   <=  32'b00111101110100110001000001000100 ;
        1098:  q   <=  32'b00111101110100110011110000011100 ;
        1099:  q   <=  32'b00111101110100110110011111110010 ;
        1100:  q   <=  32'b00111101110100111001001111000101 ;
        1101:  q   <=  32'b00111101110100111011111110010110 ;
        1102:  q   <=  32'b00111101110100111110101101100101 ;
        1103:  q   <=  32'b00111101110101000001011100110010 ;
        1104:  q   <=  32'b00111101110101000100001011111101 ;
        1105:  q   <=  32'b00111101110101000110111011000101 ;
        1106:  q   <=  32'b00111101110101001001101010001100 ;
        1107:  q   <=  32'b00111101110101001100011001010000 ;
        1108:  q   <=  32'b00111101110101001111001000010010 ;
        1109:  q   <=  32'b00111101110101010001110111010010 ;
        1110:  q   <=  32'b00111101110101010100100110010000 ;
        1111:  q   <=  32'b00111101110101010111010101001011 ;
        1112:  q   <=  32'b00111101110101011010000100000101 ;
        1113:  q   <=  32'b00111101110101011100110010111100 ;
        1114:  q   <=  32'b00111101110101011111100001110001 ;
        1115:  q   <=  32'b00111101110101100010010000100100 ;
        1116:  q   <=  32'b00111101110101100100111111010101 ;
        1117:  q   <=  32'b00111101110101100111101110000100 ;
        1118:  q   <=  32'b00111101110101101010011100110000 ;
        1119:  q   <=  32'b00111101110101101101001011011011 ;
        1120:  q   <=  32'b00111101110101101111111010000011 ;
        1121:  q   <=  32'b00111101110101110010101000101001 ;
        1122:  q   <=  32'b00111101110101110101010111001101 ;
        1123:  q   <=  32'b00111101110101111000000101101111 ;
        1124:  q   <=  32'b00111101110101111010110100001111 ;
        1125:  q   <=  32'b00111101110101111101100010101101 ;
        1126:  q   <=  32'b00111101110110000000010001001000 ;
        1127:  q   <=  32'b00111101110110000010111111100001 ;
        1128:  q   <=  32'b00111101110110000101101101111001 ;
        1129:  q   <=  32'b00111101110110001000011100001110 ;
        1130:  q   <=  32'b00111101110110001011001010100000 ;
        1131:  q   <=  32'b00111101110110001101111000110001 ;
        1132:  q   <=  32'b00111101110110010000100111000000 ;
        1133:  q   <=  32'b00111101110110010011010101001100 ;
        1134:  q   <=  32'b00111101110110010110000011010111 ;
        1135:  q   <=  32'b00111101110110011000110001011111 ;
        1136:  q   <=  32'b00111101110110011011011111100101 ;
        1137:  q   <=  32'b00111101110110011110001101101001 ;
        1138:  q   <=  32'b00111101110110100000111011101011 ;
        1139:  q   <=  32'b00111101110110100011101001101011 ;
        1140:  q   <=  32'b00111101110110100110010111101000 ;
        1141:  q   <=  32'b00111101110110101001000101100100 ;
        1142:  q   <=  32'b00111101110110101011110011011101 ;
        1143:  q   <=  32'b00111101110110101110100001010100 ;
        1144:  q   <=  32'b00111101110110110001001111001010 ;
        1145:  q   <=  32'b00111101110110110011111100111101 ;
        1146:  q   <=  32'b00111101110110110110101010101101 ;
        1147:  q   <=  32'b00111101110110111001011000011100 ;
        1148:  q   <=  32'b00111101110110111100000110001001 ;
        1149:  q   <=  32'b00111101110110111110110011110011 ;
        1150:  q   <=  32'b00111101110111000001100001011100 ;
        1151:  q   <=  32'b00111101110111000100001111000010 ;
        1152:  q   <=  32'b00111101110111000110111100100110 ;
        1153:  q   <=  32'b00111101110111001001101010001000 ;
        1154:  q   <=  32'b00111101110111001100010111101000 ;
        1155:  q   <=  32'b00111101110111001111000101000110 ;
        1156:  q   <=  32'b00111101110111010001110010100010 ;
        1157:  q   <=  32'b00111101110111010100011111111011 ;
        1158:  q   <=  32'b00111101110111010111001101010011 ;
        1159:  q   <=  32'b00111101110111011001111010101000 ;
        1160:  q   <=  32'b00111101110111011100100111111011 ;
        1161:  q   <=  32'b00111101110111011111010101001100 ;
        1162:  q   <=  32'b00111101110111100010000010011011 ;
        1163:  q   <=  32'b00111101110111100100101111101000 ;
        1164:  q   <=  32'b00111101110111100111011100110011 ;
        1165:  q   <=  32'b00111101110111101010001001111100 ;
        1166:  q   <=  32'b00111101110111101100110111000010 ;
        1167:  q   <=  32'b00111101110111101111100100000111 ;
        1168:  q   <=  32'b00111101110111110010010001001001 ;
        1169:  q   <=  32'b00111101110111110100111110001010 ;
        1170:  q   <=  32'b00111101110111110111101011001000 ;
        1171:  q   <=  32'b00111101110111111010011000000100 ;
        1172:  q   <=  32'b00111101110111111101000100111110 ;
        1173:  q   <=  32'b00111101110111111111110001110110 ;
        1174:  q   <=  32'b00111101111000000010011110101011 ;
        1175:  q   <=  32'b00111101111000000101001011011111 ;
        1176:  q   <=  32'b00111101111000000111111000010001 ;
        1177:  q   <=  32'b00111101111000001010100101000000 ;
        1178:  q   <=  32'b00111101111000001101010001101110 ;
        1179:  q   <=  32'b00111101111000001111111110011001 ;
        1180:  q   <=  32'b00111101111000010010101011000010 ;
        1181:  q   <=  32'b00111101111000010101010111101001 ;
        1182:  q   <=  32'b00111101111000011000000100001110 ;
        1183:  q   <=  32'b00111101111000011010110000110001 ;
        1184:  q   <=  32'b00111101111000011101011101010010 ;
        1185:  q   <=  32'b00111101111000100000001001110001 ;
        1186:  q   <=  32'b00111101111000100010110110001101 ;
        1187:  q   <=  32'b00111101111000100101100010101000 ;
        1188:  q   <=  32'b00111101111000101000001111000000 ;
        1189:  q   <=  32'b00111101111000101010111011010111 ;
        1190:  q   <=  32'b00111101111000101101100111101011 ;
        1191:  q   <=  32'b00111101111000110000010011111101 ;
        1192:  q   <=  32'b00111101111000110011000000001101 ;
        1193:  q   <=  32'b00111101111000110101101100011011 ;
        1194:  q   <=  32'b00111101111000111000011000100111 ;
        1195:  q   <=  32'b00111101111000111011000100110001 ;
        1196:  q   <=  32'b00111101111000111101110000111001 ;
        1197:  q   <=  32'b00111101111001000000011100111111 ;
        1198:  q   <=  32'b00111101111001000011001001000010 ;
        1199:  q   <=  32'b00111101111001000101110101000100 ;
        1200:  q   <=  32'b00111101111001001000100001000011 ;
        1201:  q   <=  32'b00111101111001001011001101000001 ;
        1202:  q   <=  32'b00111101111001001101111000111100 ;
        1203:  q   <=  32'b00111101111001010000100100110101 ;
        1204:  q   <=  32'b00111101111001010011010000101100 ;
        1205:  q   <=  32'b00111101111001010101111100100001 ;
        1206:  q   <=  32'b00111101111001011000101000010100 ;
        1207:  q   <=  32'b00111101111001011011010100000101 ;
        1208:  q   <=  32'b00111101111001011101111111110100 ;
        1209:  q   <=  32'b00111101111001100000101011100001 ;
        1210:  q   <=  32'b00111101111001100011010111001100 ;
        1211:  q   <=  32'b00111101111001100110000010110100 ;
        1212:  q   <=  32'b00111101111001101000101110011011 ;
        1213:  q   <=  32'b00111101111001101011011001111111 ;
        1214:  q   <=  32'b00111101111001101110000101100010 ;
        1215:  q   <=  32'b00111101111001110000110001000010 ;
        1216:  q   <=  32'b00111101111001110011011100100000 ;
        1217:  q   <=  32'b00111101111001110110000111111101 ;
        1218:  q   <=  32'b00111101111001111000110011010111 ;
        1219:  q   <=  32'b00111101111001111011011110101111 ;
        1220:  q   <=  32'b00111101111001111110001010000101 ;
        1221:  q   <=  32'b00111101111010000000110101011001 ;
        1222:  q   <=  32'b00111101111010000011100000101011 ;
        1223:  q   <=  32'b00111101111010000110001011111011 ;
        1224:  q   <=  32'b00111101111010001000110111001001 ;
        1225:  q   <=  32'b00111101111010001011100010010100 ;
        1226:  q   <=  32'b00111101111010001110001101011110 ;
        1227:  q   <=  32'b00111101111010010000111000100110 ;
        1228:  q   <=  32'b00111101111010010011100011101011 ;
        1229:  q   <=  32'b00111101111010010110001110101111 ;
        1230:  q   <=  32'b00111101111010011000111001110000 ;
        1231:  q   <=  32'b00111101111010011011100100110000 ;
        1232:  q   <=  32'b00111101111010011110001111101101 ;
        1233:  q   <=  32'b00111101111010100000111010101000 ;
        1234:  q   <=  32'b00111101111010100011100101100001 ;
        1235:  q   <=  32'b00111101111010100110010000011001 ;
        1236:  q   <=  32'b00111101111010101000111011001110 ;
        1237:  q   <=  32'b00111101111010101011100110000001 ;
        1238:  q   <=  32'b00111101111010101110010000110010 ;
        1239:  q   <=  32'b00111101111010110000111011100001 ;
        1240:  q   <=  32'b00111101111010110011100110001110 ;
        1241:  q   <=  32'b00111101111010110110010000111001 ;
        1242:  q   <=  32'b00111101111010111000111011100010 ;
        1243:  q   <=  32'b00111101111010111011100110001000 ;
        1244:  q   <=  32'b00111101111010111110010000101101 ;
        1245:  q   <=  32'b00111101111011000000111011010000 ;
        1246:  q   <=  32'b00111101111011000011100101110000 ;
        1247:  q   <=  32'b00111101111011000110010000001111 ;
        1248:  q   <=  32'b00111101111011001000111010101100 ;
        1249:  q   <=  32'b00111101111011001011100101000110 ;
        1250:  q   <=  32'b00111101111011001110001111011111 ;
        1251:  q   <=  32'b00111101111011010000111001110101 ;
        1252:  q   <=  32'b00111101111011010011100100001010 ;
        1253:  q   <=  32'b00111101111011010110001110011100 ;
        1254:  q   <=  32'b00111101111011011000111000101100 ;
        1255:  q   <=  32'b00111101111011011011100010111011 ;
        1256:  q   <=  32'b00111101111011011110001101000111 ;
        1257:  q   <=  32'b00111101111011100000110111010001 ;
        1258:  q   <=  32'b00111101111011100011100001011001 ;
        1259:  q   <=  32'b00111101111011100110001011100000 ;
        1260:  q   <=  32'b00111101111011101000110101100100 ;
        1261:  q   <=  32'b00111101111011101011011111100110 ;
        1262:  q   <=  32'b00111101111011101110001001100110 ;
        1263:  q   <=  32'b00111101111011110000110011100100 ;
        1264:  q   <=  32'b00111101111011110011011101100000 ;
        1265:  q   <=  32'b00111101111011110110000111011010 ;
        1266:  q   <=  32'b00111101111011111000110001010010 ;
        1267:  q   <=  32'b00111101111011111011011011001000 ;
        1268:  q   <=  32'b00111101111011111110000100111100 ;
        1269:  q   <=  32'b00111101111100000000101110101110 ;
        1270:  q   <=  32'b00111101111100000011011000011110 ;
        1271:  q   <=  32'b00111101111100000110000010001011 ;
        1272:  q   <=  32'b00111101111100001000101011110111 ;
        1273:  q   <=  32'b00111101111100001011010101100001 ;
        1274:  q   <=  32'b00111101111100001101111111001001 ;
        1275:  q   <=  32'b00111101111100010000101000101110 ;
        1276:  q   <=  32'b00111101111100010011010010010010 ;
        1277:  q   <=  32'b00111101111100010101111011110100 ;
        1278:  q   <=  32'b00111101111100011000100101010100 ;
        1279:  q   <=  32'b00111101111100011011001110110001 ;
        1280:  q   <=  32'b00111101111100011101111000001101 ;
        1281:  q   <=  32'b00111101111100100000100001100110 ;
        1282:  q   <=  32'b00111101111100100011001010111110 ;
        1283:  q   <=  32'b00111101111100100101110100010100 ;
        1284:  q   <=  32'b00111101111100101000011101100111 ;
        1285:  q   <=  32'b00111101111100101011000110111001 ;
        1286:  q   <=  32'b00111101111100101101110000001000 ;
        1287:  q   <=  32'b00111101111100110000011001010110 ;
        1288:  q   <=  32'b00111101111100110011000010100001 ;
        1289:  q   <=  32'b00111101111100110101101011101011 ;
        1290:  q   <=  32'b00111101111100111000010100110011 ;
        1291:  q   <=  32'b00111101111100111010111101111000 ;
        1292:  q   <=  32'b00111101111100111101100110111011 ;
        1293:  q   <=  32'b00111101111101000000001111111101 ;
        1294:  q   <=  32'b00111101111101000010111000111100 ;
        1295:  q   <=  32'b00111101111101000101100001111010 ;
        1296:  q   <=  32'b00111101111101001000001010110101 ;
        1297:  q   <=  32'b00111101111101001010110011101111 ;
        1298:  q   <=  32'b00111101111101001101011100100110 ;
        1299:  q   <=  32'b00111101111101010000000101011100 ;
        1300:  q   <=  32'b00111101111101010010101110001111 ;
        1301:  q   <=  32'b00111101111101010101010111000001 ;
        1302:  q   <=  32'b00111101111101010111111111110000 ;
        1303:  q   <=  32'b00111101111101011010101000011110 ;
        1304:  q   <=  32'b00111101111101011101010001001001 ;
        1305:  q   <=  32'b00111101111101011111111001110010 ;
        1306:  q   <=  32'b00111101111101100010100010011010 ;
        1307:  q   <=  32'b00111101111101100101001010111111 ;
        1308:  q   <=  32'b00111101111101100111110011100011 ;
        1309:  q   <=  32'b00111101111101101010011100000100 ;
        1310:  q   <=  32'b00111101111101101101000100100100 ;
        1311:  q   <=  32'b00111101111101101111101101000001 ;
        1312:  q   <=  32'b00111101111101110010010101011101 ;
        1313:  q   <=  32'b00111101111101110100111101110110 ;
        1314:  q   <=  32'b00111101111101110111100110001110 ;
        1315:  q   <=  32'b00111101111101111010001110100011 ;
        1316:  q   <=  32'b00111101111101111100110110110111 ;
        1317:  q   <=  32'b00111101111101111111011111001000 ;
        1318:  q   <=  32'b00111101111110000010000111011000 ;
        1319:  q   <=  32'b00111101111110000100101111100101 ;
        1320:  q   <=  32'b00111101111110000111010111110001 ;
        1321:  q   <=  32'b00111101111110001001111111111010 ;
        1322:  q   <=  32'b00111101111110001100101000000010 ;
        1323:  q   <=  32'b00111101111110001111010000001000 ;
        1324:  q   <=  32'b00111101111110010001111000001011 ;
        1325:  q   <=  32'b00111101111110010100100000001101 ;
        1326:  q   <=  32'b00111101111110010111001000001100 ;
        1327:  q   <=  32'b00111101111110011001110000001010 ;
        1328:  q   <=  32'b00111101111110011100011000000110 ;
        1329:  q   <=  32'b00111101111110011110111111111111 ;
        1330:  q   <=  32'b00111101111110100001100111110111 ;
        1331:  q   <=  32'b00111101111110100100001111101101 ;
        1332:  q   <=  32'b00111101111110100110110111100001 ;
        1333:  q   <=  32'b00111101111110101001011111010010 ;
        1334:  q   <=  32'b00111101111110101100000111000010 ;
        1335:  q   <=  32'b00111101111110101110101110110000 ;
        1336:  q   <=  32'b00111101111110110001010110011100 ;
        1337:  q   <=  32'b00111101111110110011111110000110 ;
        1338:  q   <=  32'b00111101111110110110100101101110 ;
        1339:  q   <=  32'b00111101111110111001001101010100 ;
        1340:  q   <=  32'b00111101111110111011110100111000 ;
        1341:  q   <=  32'b00111101111110111110011100011010 ;
        1342:  q   <=  32'b00111101111111000001000011111010 ;
        1343:  q   <=  32'b00111101111111000011101011011000 ;
        1344:  q   <=  32'b00111101111111000110010010110100 ;
        1345:  q   <=  32'b00111101111111001000111010001110 ;
        1346:  q   <=  32'b00111101111111001011100001100110 ;
        1347:  q   <=  32'b00111101111111001110001000111100 ;
        1348:  q   <=  32'b00111101111111010000110000010000 ;
        1349:  q   <=  32'b00111101111111010011010111100010 ;
        1350:  q   <=  32'b00111101111111010101111110110011 ;
        1351:  q   <=  32'b00111101111111011000100110000001 ;
        1352:  q   <=  32'b00111101111111011011001101001101 ;
        1353:  q   <=  32'b00111101111111011101110100011000 ;
        1354:  q   <=  32'b00111101111111100000011011100000 ;
        1355:  q   <=  32'b00111101111111100011000010100110 ;
        1356:  q   <=  32'b00111101111111100101101001101011 ;
        1357:  q   <=  32'b00111101111111101000010000101101 ;
        1358:  q   <=  32'b00111101111111101010110111101110 ;
        1359:  q   <=  32'b00111101111111101101011110101101 ;
        1360:  q   <=  32'b00111101111111110000000101101001 ;
        1361:  q   <=  32'b00111101111111110010101100100100 ;
        1362:  q   <=  32'b00111101111111110101010011011101 ;
        1363:  q   <=  32'b00111101111111110111111010010011 ;
        1364:  q   <=  32'b00111101111111111010100001001000 ;
        1365:  q   <=  32'b00111101111111111101000111111011 ;
        1366:  q   <=  32'b00111101111111111111101110101100 ;
        1367:  q   <=  32'b00111110000000000001001010101101 ;
        1368:  q   <=  32'b00111110000000000010011110000100 ;
        1369:  q   <=  32'b00111110000000000011110001011001 ;
        1370:  q   <=  32'b00111110000000000101000100101110 ;
        1371:  q   <=  32'b00111110000000000110011000000001 ;
        1372:  q   <=  32'b00111110000000000111101011010100 ;
        1373:  q   <=  32'b00111110000000001000111110100110 ;
        1374:  q   <=  32'b00111110000000001010010001110110 ;
        1375:  q   <=  32'b00111110000000001011100101000110 ;
        1376:  q   <=  32'b00111110000000001100111000010101 ;
        1377:  q   <=  32'b00111110000000001110001011100010 ;
        1378:  q   <=  32'b00111110000000001111011110101111 ;
        1379:  q   <=  32'b00111110000000010000110001111011 ;
        1380:  q   <=  32'b00111110000000010010000101000110 ;
        1381:  q   <=  32'b00111110000000010011011000001111 ;
        1382:  q   <=  32'b00111110000000010100101011011000 ;
        1383:  q   <=  32'b00111110000000010101111110100000 ;
        1384:  q   <=  32'b00111110000000010111010001100111 ;
        1385:  q   <=  32'b00111110000000011000100100101101 ;
        1386:  q   <=  32'b00111110000000011001110111110010 ;
        1387:  q   <=  32'b00111110000000011011001010110110 ;
        1388:  q   <=  32'b00111110000000011100011101111001 ;
        1389:  q   <=  32'b00111110000000011101110000111011 ;
        1390:  q   <=  32'b00111110000000011111000011111100 ;
        1391:  q   <=  32'b00111110000000100000010110111100 ;
        1392:  q   <=  32'b00111110000000100001101001111011 ;
        1393:  q   <=  32'b00111110000000100010111100111010 ;
        1394:  q   <=  32'b00111110000000100100001111110111 ;
        1395:  q   <=  32'b00111110000000100101100010110011 ;
        1396:  q   <=  32'b00111110000000100110110101101110 ;
        1397:  q   <=  32'b00111110000000101000001000101001 ;
        1398:  q   <=  32'b00111110000000101001011011100010 ;
        1399:  q   <=  32'b00111110000000101010101110011011 ;
        1400:  q   <=  32'b00111110000000101100000001010010 ;
        1401:  q   <=  32'b00111110000000101101010100001000 ;
        1402:  q   <=  32'b00111110000000101110100110111110 ;
        1403:  q   <=  32'b00111110000000101111111001110010 ;
        1404:  q   <=  32'b00111110000000110001001100100110 ;
        1405:  q   <=  32'b00111110000000110010011111011001 ;
        1406:  q   <=  32'b00111110000000110011110010001010 ;
        1407:  q   <=  32'b00111110000000110101000100111011 ;
        1408:  q   <=  32'b00111110000000110110010111101011 ;
        1409:  q   <=  32'b00111110000000110111101010011001 ;
        1410:  q   <=  32'b00111110000000111000111101000111 ;
        1411:  q   <=  32'b00111110000000111010001111110100 ;
        1412:  q   <=  32'b00111110000000111011100010100000 ;
        1413:  q   <=  32'b00111110000000111100110101001011 ;
        1414:  q   <=  32'b00111110000000111110000111110101 ;
        1415:  q   <=  32'b00111110000000111111011010011110 ;
        1416:  q   <=  32'b00111110000001000000101101000110 ;
        1417:  q   <=  32'b00111110000001000001111111101101 ;
        1418:  q   <=  32'b00111110000001000011010010010011 ;
        1419:  q   <=  32'b00111110000001000100100100111000 ;
        1420:  q   <=  32'b00111110000001000101110111011100 ;
        1421:  q   <=  32'b00111110000001000111001010000000 ;
        1422:  q   <=  32'b00111110000001001000011100100010 ;
        1423:  q   <=  32'b00111110000001001001101111000011 ;
        1424:  q   <=  32'b00111110000001001011000001100100 ;
        1425:  q   <=  32'b00111110000001001100010100000011 ;
        1426:  q   <=  32'b00111110000001001101100110100010 ;
        1427:  q   <=  32'b00111110000001001110111000111111 ;
        1428:  q   <=  32'b00111110000001010000001011011100 ;
        1429:  q   <=  32'b00111110000001010001011101110111 ;
        1430:  q   <=  32'b00111110000001010010110000010010 ;
        1431:  q   <=  32'b00111110000001010100000010101100 ;
        1432:  q   <=  32'b00111110000001010101010101000100 ;
        1433:  q   <=  32'b00111110000001010110100111011100 ;
        1434:  q   <=  32'b00111110000001010111111001110011 ;
        1435:  q   <=  32'b00111110000001011001001100001001 ;
        1436:  q   <=  32'b00111110000001011010011110011110 ;
        1437:  q   <=  32'b00111110000001011011110000110010 ;
        1438:  q   <=  32'b00111110000001011101000011000101 ;
        1439:  q   <=  32'b00111110000001011110010101010111 ;
        1440:  q   <=  32'b00111110000001011111100111101000 ;
        1441:  q   <=  32'b00111110000001100000111001111000 ;
        1442:  q   <=  32'b00111110000001100010001100000111 ;
        1443:  q   <=  32'b00111110000001100011011110010101 ;
        1444:  q   <=  32'b00111110000001100100110000100011 ;
        1445:  q   <=  32'b00111110000001100110000010101111 ;
        1446:  q   <=  32'b00111110000001100111010100111010 ;
        1447:  q   <=  32'b00111110000001101000100111000101 ;
        1448:  q   <=  32'b00111110000001101001111001001110 ;
        1449:  q   <=  32'b00111110000001101011001011010111 ;
        1450:  q   <=  32'b00111110000001101100011101011111 ;
        1451:  q   <=  32'b00111110000001101101101111100101 ;
        1452:  q   <=  32'b00111110000001101111000001101011 ;
        1453:  q   <=  32'b00111110000001110000010011110000 ;
        1454:  q   <=  32'b00111110000001110001100101110100 ;
        1455:  q   <=  32'b00111110000001110010110111110110 ;
        1456:  q   <=  32'b00111110000001110100001001111000 ;
        1457:  q   <=  32'b00111110000001110101011011111001 ;
        1458:  q   <=  32'b00111110000001110110101101111001 ;
        1459:  q   <=  32'b00111110000001110111111111111001 ;
        1460:  q   <=  32'b00111110000001111001010001110111 ;
        1461:  q   <=  32'b00111110000001111010100011110100 ;
        1462:  q   <=  32'b00111110000001111011110101110000 ;
        1463:  q   <=  32'b00111110000001111101000111101100 ;
        1464:  q   <=  32'b00111110000001111110011001100110 ;
        1465:  q   <=  32'b00111110000001111111101011011111 ;
        1466:  q   <=  32'b00111110000010000000111101011000 ;
        1467:  q   <=  32'b00111110000010000010001111001111 ;
        1468:  q   <=  32'b00111110000010000011100001000110 ;
        1469:  q   <=  32'b00111110000010000100110010111100 ;
        1470:  q   <=  32'b00111110000010000110000100110000 ;
        1471:  q   <=  32'b00111110000010000111010110100100 ;
        1472:  q   <=  32'b00111110000010001000101000010111 ;
        1473:  q   <=  32'b00111110000010001001111010001001 ;
        1474:  q   <=  32'b00111110000010001011001011111010 ;
        1475:  q   <=  32'b00111110000010001100011101101010 ;
        1476:  q   <=  32'b00111110000010001101101111011001 ;
        1477:  q   <=  32'b00111110000010001111000001000111 ;
        1478:  q   <=  32'b00111110000010010000010010110100 ;
        1479:  q   <=  32'b00111110000010010001100100100001 ;
        1480:  q   <=  32'b00111110000010010010110110001100 ;
        1481:  q   <=  32'b00111110000010010100000111110110 ;
        1482:  q   <=  32'b00111110000010010101011001100000 ;
        1483:  q   <=  32'b00111110000010010110101011001000 ;
        1484:  q   <=  32'b00111110000010010111111100110000 ;
        1485:  q   <=  32'b00111110000010011001001110010111 ;
        1486:  q   <=  32'b00111110000010011010011111111100 ;
        1487:  q   <=  32'b00111110000010011011110001100001 ;
        1488:  q   <=  32'b00111110000010011101000011000101 ;
        1489:  q   <=  32'b00111110000010011110010100101000 ;
        1490:  q   <=  32'b00111110000010011111100110001010 ;
        1491:  q   <=  32'b00111110000010100000110111101011 ;
        1492:  q   <=  32'b00111110000010100010001001001011 ;
        1493:  q   <=  32'b00111110000010100011011010101010 ;
        1494:  q   <=  32'b00111110000010100100101100001000 ;
        1495:  q   <=  32'b00111110000010100101111101100110 ;
        1496:  q   <=  32'b00111110000010100111001111000010 ;
        1497:  q   <=  32'b00111110000010101000100000011110 ;
        1498:  q   <=  32'b00111110000010101001110001111000 ;
        1499:  q   <=  32'b00111110000010101011000011010010 ;
        1500:  q   <=  32'b00111110000010101100010100101010 ;
        1501:  q   <=  32'b00111110000010101101100110000010 ;
        1502:  q   <=  32'b00111110000010101110110111011001 ;
        1503:  q   <=  32'b00111110000010110000001000101111 ;
        1504:  q   <=  32'b00111110000010110001011010000100 ;
        1505:  q   <=  32'b00111110000010110010101011011000 ;
        1506:  q   <=  32'b00111110000010110011111100101011 ;
        1507:  q   <=  32'b00111110000010110101001101111101 ;
        1508:  q   <=  32'b00111110000010110110011111001110 ;
        1509:  q   <=  32'b00111110000010110111110000011110 ;
        1510:  q   <=  32'b00111110000010111001000001101110 ;
        1511:  q   <=  32'b00111110000010111010010010111100 ;
        1512:  q   <=  32'b00111110000010111011100100001010 ;
        1513:  q   <=  32'b00111110000010111100110101010110 ;
        1514:  q   <=  32'b00111110000010111110000110100010 ;
        1515:  q   <=  32'b00111110000010111111010111101101 ;
        1516:  q   <=  32'b00111110000011000000101000110110 ;
        1517:  q   <=  32'b00111110000011000001111001111111 ;
        1518:  q   <=  32'b00111110000011000011001011000111 ;
        1519:  q   <=  32'b00111110000011000100011100001110 ;
        1520:  q   <=  32'b00111110000011000101101101010100 ;
        1521:  q   <=  32'b00111110000011000110111110011001 ;
        1522:  q   <=  32'b00111110000011001000001111011110 ;
        1523:  q   <=  32'b00111110000011001001100000100001 ;
        1524:  q   <=  32'b00111110000011001010110001100011 ;
        1525:  q   <=  32'b00111110000011001100000010100101 ;
        1526:  q   <=  32'b00111110000011001101010011100110 ;
        1527:  q   <=  32'b00111110000011001110100100100101 ;
        1528:  q   <=  32'b00111110000011001111110101100100 ;
        1529:  q   <=  32'b00111110000011010001000110100010 ;
        1530:  q   <=  32'b00111110000011010010010111011111 ;
        1531:  q   <=  32'b00111110000011010011101000011010 ;
        1532:  q   <=  32'b00111110000011010100111001010110 ;
        1533:  q   <=  32'b00111110000011010110001010010000 ;
        1534:  q   <=  32'b00111110000011010111011011001001 ;
        1535:  q   <=  32'b00111110000011011000101100000001 ;
        1536:  q   <=  32'b00111110000011011001111100111000 ;
        1537:  q   <=  32'b00111110000011011011001101101111 ;
        1538:  q   <=  32'b00111110000011011100011110100100 ;
        1539:  q   <=  32'b00111110000011011101101111011001 ;
        1540:  q   <=  32'b00111110000011011111000000001101 ;
        1541:  q   <=  32'b00111110000011100000010000111111 ;
        1542:  q   <=  32'b00111110000011100001100001110001 ;
        1543:  q   <=  32'b00111110000011100010110010100010 ;
        1544:  q   <=  32'b00111110000011100100000011010010 ;
        1545:  q   <=  32'b00111110000011100101010100000001 ;
        1546:  q   <=  32'b00111110000011100110100100110000 ;
        1547:  q   <=  32'b00111110000011100111110101011101 ;
        1548:  q   <=  32'b00111110000011101001000110001001 ;
        1549:  q   <=  32'b00111110000011101010010110110101 ;
        1550:  q   <=  32'b00111110000011101011100111011111 ;
        1551:  q   <=  32'b00111110000011101100111000001001 ;
        1552:  q   <=  32'b00111110000011101110001000110001 ;
        1553:  q   <=  32'b00111110000011101111011001011001 ;
        1554:  q   <=  32'b00111110000011110000101010000000 ;
        1555:  q   <=  32'b00111110000011110001111010100110 ;
        1556:  q   <=  32'b00111110000011110011001011001011 ;
        1557:  q   <=  32'b00111110000011110100011011101111 ;
        1558:  q   <=  32'b00111110000011110101101100010010 ;
        1559:  q   <=  32'b00111110000011110110111100110101 ;
        1560:  q   <=  32'b00111110000011111000001101010110 ;
        1561:  q   <=  32'b00111110000011111001011101110111 ;
        1562:  q   <=  32'b00111110000011111010101110010110 ;
        1563:  q   <=  32'b00111110000011111011111110110101 ;
        1564:  q   <=  32'b00111110000011111101001111010011 ;
        1565:  q   <=  32'b00111110000011111110011111101111 ;
        1566:  q   <=  32'b00111110000011111111110000001011 ;
        1567:  q   <=  32'b00111110000100000001000000100110 ;
        1568:  q   <=  32'b00111110000100000010010001000000 ;
        1569:  q   <=  32'b00111110000100000011100001011010 ;
        1570:  q   <=  32'b00111110000100000100110001110010 ;
        1571:  q   <=  32'b00111110000100000110000010001001 ;
        1572:  q   <=  32'b00111110000100000111010010100000 ;
        1573:  q   <=  32'b00111110000100001000100010110101 ;
        1574:  q   <=  32'b00111110000100001001110011001010 ;
        1575:  q   <=  32'b00111110000100001011000011011110 ;
        1576:  q   <=  32'b00111110000100001100010011110001 ;
        1577:  q   <=  32'b00111110000100001101100100000011 ;
        1578:  q   <=  32'b00111110000100001110110100010100 ;
        1579:  q   <=  32'b00111110000100010000000100100100 ;
        1580:  q   <=  32'b00111110000100010001010100110011 ;
        1581:  q   <=  32'b00111110000100010010100101000001 ;
        1582:  q   <=  32'b00111110000100010011110101001111 ;
        1583:  q   <=  32'b00111110000100010101000101011011 ;
        1584:  q   <=  32'b00111110000100010110010101100111 ;
        1585:  q   <=  32'b00111110000100010111100101110010 ;
        1586:  q   <=  32'b00111110000100011000110101111011 ;
        1587:  q   <=  32'b00111110000100011010000110000100 ;
        1588:  q   <=  32'b00111110000100011011010110001100 ;
        1589:  q   <=  32'b00111110000100011100100110010011 ;
        1590:  q   <=  32'b00111110000100011101110110011010 ;
        1591:  q   <=  32'b00111110000100011111000110011111 ;
        1592:  q   <=  32'b00111110000100100000010110100011 ;
        1593:  q   <=  32'b00111110000100100001100110100111 ;
        1594:  q   <=  32'b00111110000100100010110110101001 ;
        1595:  q   <=  32'b00111110000100100100000110101011 ;
        1596:  q   <=  32'b00111110000100100101010110101100 ;
        1597:  q   <=  32'b00111110000100100110100110101100 ;
        1598:  q   <=  32'b00111110000100100111110110101011 ;
        1599:  q   <=  32'b00111110000100101001000110101001 ;
        1600:  q   <=  32'b00111110000100101010010110100110 ;
        1601:  q   <=  32'b00111110000100101011100110100010 ;
        1602:  q   <=  32'b00111110000100101100110110011110 ;
        1603:  q   <=  32'b00111110000100101110000110011000 ;
        1604:  q   <=  32'b00111110000100101111010110010010 ;
        1605:  q   <=  32'b00111110000100110000100110001011 ;
        1606:  q   <=  32'b00111110000100110001110110000010 ;
        1607:  q   <=  32'b00111110000100110011000101111001 ;
        1608:  q   <=  32'b00111110000100110100010101101111 ;
        1609:  q   <=  32'b00111110000100110101100101100101 ;
        1610:  q   <=  32'b00111110000100110110110101011001 ;
        1611:  q   <=  32'b00111110000100111000000101001100 ;
        1612:  q   <=  32'b00111110000100111001010100111111 ;
        1613:  q   <=  32'b00111110000100111010100100110000 ;
        1614:  q   <=  32'b00111110000100111011110100100001 ;
        1615:  q   <=  32'b00111110000100111101000100010000 ;
        1616:  q   <=  32'b00111110000100111110010011111111 ;
        1617:  q   <=  32'b00111110000100111111100011101101 ;
        1618:  q   <=  32'b00111110000101000000110011011010 ;
        1619:  q   <=  32'b00111110000101000010000011000111 ;
        1620:  q   <=  32'b00111110000101000011010010110010 ;
        1621:  q   <=  32'b00111110000101000100100010011100 ;
        1622:  q   <=  32'b00111110000101000101110010000110 ;
        1623:  q   <=  32'b00111110000101000111000001101110 ;
        1624:  q   <=  32'b00111110000101001000010001010110 ;
        1625:  q   <=  32'b00111110000101001001100000111101 ;
        1626:  q   <=  32'b00111110000101001010110000100011 ;
        1627:  q   <=  32'b00111110000101001100000000001000 ;
        1628:  q   <=  32'b00111110000101001101001111101100 ;
        1629:  q   <=  32'b00111110000101001110011111001111 ;
        1630:  q   <=  32'b00111110000101001111101110110010 ;
        1631:  q   <=  32'b00111110000101010000111110010011 ;
        1632:  q   <=  32'b00111110000101010010001101110100 ;
        1633:  q   <=  32'b00111110000101010011011101010100 ;
        1634:  q   <=  32'b00111110000101010100101100110010 ;
        1635:  q   <=  32'b00111110000101010101111100010000 ;
        1636:  q   <=  32'b00111110000101010111001011101101 ;
        1637:  q   <=  32'b00111110000101011000011011001010 ;
        1638:  q   <=  32'b00111110000101011001101010100101 ;
        1639:  q   <=  32'b00111110000101011010111001111111 ;
        1640:  q   <=  32'b00111110000101011100001001011001 ;
        1641:  q   <=  32'b00111110000101011101011000110001 ;
        1642:  q   <=  32'b00111110000101011110101000001001 ;
        1643:  q   <=  32'b00111110000101011111110111100000 ;
        1644:  q   <=  32'b00111110000101100001000110110110 ;
        1645:  q   <=  32'b00111110000101100010010110001011 ;
        1646:  q   <=  32'b00111110000101100011100101011111 ;
        1647:  q   <=  32'b00111110000101100100110100110011 ;
        1648:  q   <=  32'b00111110000101100110000100000101 ;
        1649:  q   <=  32'b00111110000101100111010011010111 ;
        1650:  q   <=  32'b00111110000101101000100010100111 ;
        1651:  q   <=  32'b00111110000101101001110001110111 ;
        1652:  q   <=  32'b00111110000101101011000001000110 ;
        1653:  q   <=  32'b00111110000101101100010000010100 ;
        1654:  q   <=  32'b00111110000101101101011111100001 ;
        1655:  q   <=  32'b00111110000101101110101110101101 ;
        1656:  q   <=  32'b00111110000101101111111101111001 ;
        1657:  q   <=  32'b00111110000101110001001101000011 ;
        1658:  q   <=  32'b00111110000101110010011100001101 ;
        1659:  q   <=  32'b00111110000101110011101011010110 ;
        1660:  q   <=  32'b00111110000101110100111010011101 ;
        1661:  q   <=  32'b00111110000101110110001001100100 ;
        1662:  q   <=  32'b00111110000101110111011000101011 ;
        1663:  q   <=  32'b00111110000101111000100111110000 ;
        1664:  q   <=  32'b00111110000101111001110110110100 ;
        1665:  q   <=  32'b00111110000101111011000101111000 ;
        1666:  q   <=  32'b00111110000101111100010100111010 ;
        1667:  q   <=  32'b00111110000101111101100011111100 ;
        1668:  q   <=  32'b00111110000101111110110010111101 ;
        1669:  q   <=  32'b00111110000110000000000001111101 ;
        1670:  q   <=  32'b00111110000110000001010000111100 ;
        1671:  q   <=  32'b00111110000110000010011111111010 ;
        1672:  q   <=  32'b00111110000110000011101110110111 ;
        1673:  q   <=  32'b00111110000110000100111101110100 ;
        1674:  q   <=  32'b00111110000110000110001100101111 ;
        1675:  q   <=  32'b00111110000110000111011011101010 ;
        1676:  q   <=  32'b00111110000110001000101010100100 ;
        1677:  q   <=  32'b00111110000110001001111001011101 ;
        1678:  q   <=  32'b00111110000110001011001000010101 ;
        1679:  q   <=  32'b00111110000110001100010111001100 ;
        1680:  q   <=  32'b00111110000110001101100110000010 ;
        1681:  q   <=  32'b00111110000110001110110100111000 ;
        1682:  q   <=  32'b00111110000110010000000011101100 ;
        1683:  q   <=  32'b00111110000110010001010010100000 ;
        1684:  q   <=  32'b00111110000110010010100001010011 ;
        1685:  q   <=  32'b00111110000110010011110000000101 ;
        1686:  q   <=  32'b00111110000110010100111110110110 ;
        1687:  q   <=  32'b00111110000110010110001101100110 ;
        1688:  q   <=  32'b00111110000110010111011100010101 ;
        1689:  q   <=  32'b00111110000110011000101011000100 ;
        1690:  q   <=  32'b00111110000110011001111001110001 ;
        1691:  q   <=  32'b00111110000110011011001000011110 ;
        1692:  q   <=  32'b00111110000110011100010111001010 ;
        1693:  q   <=  32'b00111110000110011101100101110101 ;
        1694:  q   <=  32'b00111110000110011110110100011111 ;
        1695:  q   <=  32'b00111110000110100000000011001000 ;
        1696:  q   <=  32'b00111110000110100001010001110001 ;
        1697:  q   <=  32'b00111110000110100010100000011000 ;
        1698:  q   <=  32'b00111110000110100011101110111111 ;
        1699:  q   <=  32'b00111110000110100100111101100101 ;
        1700:  q   <=  32'b00111110000110100110001100001001 ;
        1701:  q   <=  32'b00111110000110100111011010101110 ;
        1702:  q   <=  32'b00111110000110101000101001010001 ;
        1703:  q   <=  32'b00111110000110101001110111110011 ;
        1704:  q   <=  32'b00111110000110101011000110010100 ;
        1705:  q   <=  32'b00111110000110101100010100110101 ;
        1706:  q   <=  32'b00111110000110101101100011010101 ;
        1707:  q   <=  32'b00111110000110101110110001110100 ;
        1708:  q   <=  32'b00111110000110110000000000010010 ;
        1709:  q   <=  32'b00111110000110110001001110101111 ;
        1710:  q   <=  32'b00111110000110110010011101001011 ;
        1711:  q   <=  32'b00111110000110110011101011100110 ;
        1712:  q   <=  32'b00111110000110110100111010000001 ;
        1713:  q   <=  32'b00111110000110110110001000011010 ;
        1714:  q   <=  32'b00111110000110110111010110110011 ;
        1715:  q   <=  32'b00111110000110111000100101001011 ;
        1716:  q   <=  32'b00111110000110111001110011100010 ;
        1717:  q   <=  32'b00111110000110111011000001111000 ;
        1718:  q   <=  32'b00111110000110111100010000001110 ;
        1719:  q   <=  32'b00111110000110111101011110100010 ;
        1720:  q   <=  32'b00111110000110111110101100110110 ;
        1721:  q   <=  32'b00111110000110111111111011001001 ;
        1722:  q   <=  32'b00111110000111000001001001011010 ;
        1723:  q   <=  32'b00111110000111000010010111101011 ;
        1724:  q   <=  32'b00111110000111000011100101111100 ;
        1725:  q   <=  32'b00111110000111000100110100001011 ;
        1726:  q   <=  32'b00111110000111000110000010011001 ;
        1727:  q   <=  32'b00111110000111000111010000100111 ;
        1728:  q   <=  32'b00111110000111001000011110110100 ;
        1729:  q   <=  32'b00111110000111001001101100111111 ;
        1730:  q   <=  32'b00111110000111001010111011001011 ;
        1731:  q   <=  32'b00111110000111001100001001010101 ;
        1732:  q   <=  32'b00111110000111001101010111011110 ;
        1733:  q   <=  32'b00111110000111001110100101100110 ;
        1734:  q   <=  32'b00111110000111001111110011101110 ;
        1735:  q   <=  32'b00111110000111010001000001110101 ;
        1736:  q   <=  32'b00111110000111010010001111111011 ;
        1737:  q   <=  32'b00111110000111010011011110000000 ;
        1738:  q   <=  32'b00111110000111010100101100000100 ;
        1739:  q   <=  32'b00111110000111010101111010000111 ;
        1740:  q   <=  32'b00111110000111010111001000001001 ;
        1741:  q   <=  32'b00111110000111011000010110001011 ;
        1742:  q   <=  32'b00111110000111011001100100001100 ;
        1743:  q   <=  32'b00111110000111011010110010001100 ;
        1744:  q   <=  32'b00111110000111011100000000001011 ;
        1745:  q   <=  32'b00111110000111011101001110001001 ;
        1746:  q   <=  32'b00111110000111011110011100000110 ;
        1747:  q   <=  32'b00111110000111011111101010000010 ;
        1748:  q   <=  32'b00111110000111100000110111111110 ;
        1749:  q   <=  32'b00111110000111100010000101111001 ;
        1750:  q   <=  32'b00111110000111100011010011110011 ;
        1751:  q   <=  32'b00111110000111100100100001101100 ;
        1752:  q   <=  32'b00111110000111100101101111100100 ;
        1753:  q   <=  32'b00111110000111100110111101011011 ;
        1754:  q   <=  32'b00111110000111101000001011010010 ;
        1755:  q   <=  32'b00111110000111101001011001000111 ;
        1756:  q   <=  32'b00111110000111101010100110111100 ;
        1757:  q   <=  32'b00111110000111101011110100110000 ;
        1758:  q   <=  32'b00111110000111101101000010100011 ;
        1759:  q   <=  32'b00111110000111101110010000010101 ;
        1760:  q   <=  32'b00111110000111101111011110000111 ;
        1761:  q   <=  32'b00111110000111110000101011110111 ;
        1762:  q   <=  32'b00111110000111110001111001100111 ;
        1763:  q   <=  32'b00111110000111110011000111010110 ;
        1764:  q   <=  32'b00111110000111110100010101000100 ;
        1765:  q   <=  32'b00111110000111110101100010110001 ;
        1766:  q   <=  32'b00111110000111110110110000011101 ;
        1767:  q   <=  32'b00111110000111110111111110001001 ;
        1768:  q   <=  32'b00111110000111111001001011110011 ;
        1769:  q   <=  32'b00111110000111111010011001011101 ;
        1770:  q   <=  32'b00111110000111111011100111000110 ;
        1771:  q   <=  32'b00111110000111111100110100101110 ;
        1772:  q   <=  32'b00111110000111111110000010010101 ;
        1773:  q   <=  32'b00111110000111111111001111111011 ;
        1774:  q   <=  32'b00111110001000000000011101100001 ;
        1775:  q   <=  32'b00111110001000000001101011000101 ;
        1776:  q   <=  32'b00111110001000000010111000101001 ;
        1777:  q   <=  32'b00111110001000000100000110001100 ;
        1778:  q   <=  32'b00111110001000000101010011101110 ;
        1779:  q   <=  32'b00111110001000000110100001010000 ;
        1780:  q   <=  32'b00111110001000000111101110110000 ;
        1781:  q   <=  32'b00111110001000001000111100010000 ;
        1782:  q   <=  32'b00111110001000001010001001101110 ;
        1783:  q   <=  32'b00111110001000001011010111001100 ;
        1784:  q   <=  32'b00111110001000001100100100101001 ;
        1785:  q   <=  32'b00111110001000001101110010000110 ;
        1786:  q   <=  32'b00111110001000001110111111100001 ;
        1787:  q   <=  32'b00111110001000010000001100111011 ;
        1788:  q   <=  32'b00111110001000010001011010010101 ;
        1789:  q   <=  32'b00111110001000010010100111101110 ;
        1790:  q   <=  32'b00111110001000010011110101000110 ;
        1791:  q   <=  32'b00111110001000010101000010011101 ;
        1792:  q   <=  32'b00111110001000010110001111110011 ;
        1793:  q   <=  32'b00111110001000010111011101001001 ;
        1794:  q   <=  32'b00111110001000011000101010011110 ;
        1795:  q   <=  32'b00111110001000011001110111110001 ;
        1796:  q   <=  32'b00111110001000011011000101000100 ;
        1797:  q   <=  32'b00111110001000011100010010010110 ;
        1798:  q   <=  32'b00111110001000011101011111101000 ;
        1799:  q   <=  32'b00111110001000011110101100111000 ;
        1800:  q   <=  32'b00111110001000011111111010001000 ;
        1801:  q   <=  32'b00111110001000100001000111010111 ;
        1802:  q   <=  32'b00111110001000100010010100100101 ;
        1803:  q   <=  32'b00111110001000100011100001110010 ;
        1804:  q   <=  32'b00111110001000100100101110111110 ;
        1805:  q   <=  32'b00111110001000100101111100001001 ;
        1806:  q   <=  32'b00111110001000100111001001010100 ;
        1807:  q   <=  32'b00111110001000101000010110011110 ;
        1808:  q   <=  32'b00111110001000101001100011100110 ;
        1809:  q   <=  32'b00111110001000101010110000101111 ;
        1810:  q   <=  32'b00111110001000101011111101110110 ;
        1811:  q   <=  32'b00111110001000101101001010111100 ;
        1812:  q   <=  32'b00111110001000101110011000000010 ;
        1813:  q   <=  32'b00111110001000101111100101000110 ;
        1814:  q   <=  32'b00111110001000110000110010001010 ;
        1815:  q   <=  32'b00111110001000110001111111001101 ;
        1816:  q   <=  32'b00111110001000110011001100010000 ;
        1817:  q   <=  32'b00111110001000110100011001010001 ;
        1818:  q   <=  32'b00111110001000110101100110010010 ;
        1819:  q   <=  32'b00111110001000110110110011010001 ;
        1820:  q   <=  32'b00111110001000111000000000010000 ;
        1821:  q   <=  32'b00111110001000111001001101001110 ;
        1822:  q   <=  32'b00111110001000111010011010001011 ;
        1823:  q   <=  32'b00111110001000111011100111001000 ;
        1824:  q   <=  32'b00111110001000111100110100000011 ;
        1825:  q   <=  32'b00111110001000111110000000111110 ;
        1826:  q   <=  32'b00111110001000111111001101111000 ;
        1827:  q   <=  32'b00111110001001000000011010110001 ;
        1828:  q   <=  32'b00111110001001000001100111101001 ;
        1829:  q   <=  32'b00111110001001000010110100100001 ;
        1830:  q   <=  32'b00111110001001000100000001010111 ;
        1831:  q   <=  32'b00111110001001000101001110001101 ;
        1832:  q   <=  32'b00111110001001000110011011000010 ;
        1833:  q   <=  32'b00111110001001000111100111110110 ;
        1834:  q   <=  32'b00111110001001001000110100101001 ;
        1835:  q   <=  32'b00111110001001001010000001011100 ;
        1836:  q   <=  32'b00111110001001001011001110001101 ;
        1837:  q   <=  32'b00111110001001001100011010111110 ;
        1838:  q   <=  32'b00111110001001001101100111101110 ;
        1839:  q   <=  32'b00111110001001001110110100011101 ;
        1840:  q   <=  32'b00111110001001010000000001001011 ;
        1841:  q   <=  32'b00111110001001010001001101111001 ;
        1842:  q   <=  32'b00111110001001010010011010100110 ;
        1843:  q   <=  32'b00111110001001010011100111010001 ;
        1844:  q   <=  32'b00111110001001010100110011111100 ;
        1845:  q   <=  32'b00111110001001010110000000100110 ;
        1846:  q   <=  32'b00111110001001010111001101010000 ;
        1847:  q   <=  32'b00111110001001011000011001111000 ;
        1848:  q   <=  32'b00111110001001011001100110100000 ;
        1849:  q   <=  32'b00111110001001011010110011000111 ;
        1850:  q   <=  32'b00111110001001011011111111101101 ;
        1851:  q   <=  32'b00111110001001011101001100010010 ;
        1852:  q   <=  32'b00111110001001011110011000110110 ;
        1853:  q   <=  32'b00111110001001011111100101011010 ;
        1854:  q   <=  32'b00111110001001100000110001111101 ;
        1855:  q   <=  32'b00111110001001100001111110011111 ;
        1856:  q   <=  32'b00111110001001100011001011000000 ;
        1857:  q   <=  32'b00111110001001100100010111100000 ;
        1858:  q   <=  32'b00111110001001100101100011111111 ;
        1859:  q   <=  32'b00111110001001100110110000011110 ;
        1860:  q   <=  32'b00111110001001100111111100111100 ;
        1861:  q   <=  32'b00111110001001101001001001011001 ;
        1862:  q   <=  32'b00111110001001101010010101110101 ;
        1863:  q   <=  32'b00111110001001101011100010010000 ;
        1864:  q   <=  32'b00111110001001101100101110101011 ;
        1865:  q   <=  32'b00111110001001101101111011000101 ;
        1866:  q   <=  32'b00111110001001101111000111011101 ;
        1867:  q   <=  32'b00111110001001110000010011110101 ;
        1868:  q   <=  32'b00111110001001110001100000001101 ;
        1869:  q   <=  32'b00111110001001110010101100100011 ;
        1870:  q   <=  32'b00111110001001110011111000111001 ;
        1871:  q   <=  32'b00111110001001110101000101001101 ;
        1872:  q   <=  32'b00111110001001110110010001100001 ;
        1873:  q   <=  32'b00111110001001110111011101110101 ;
        1874:  q   <=  32'b00111110001001111000101010000111 ;
        1875:  q   <=  32'b00111110001001111001110110011000 ;
        1876:  q   <=  32'b00111110001001111011000010101001 ;
        1877:  q   <=  32'b00111110001001111100001110111001 ;
        1878:  q   <=  32'b00111110001001111101011011001000 ;
        1879:  q   <=  32'b00111110001001111110100111010110 ;
        1880:  q   <=  32'b00111110001001111111110011100100 ;
        1881:  q   <=  32'b00111110001010000000111111110000 ;
        1882:  q   <=  32'b00111110001010000010001011111100 ;
        1883:  q   <=  32'b00111110001010000011011000000111 ;
        1884:  q   <=  32'b00111110001010000100100100010001 ;
        1885:  q   <=  32'b00111110001010000101110000011010 ;
        1886:  q   <=  32'b00111110001010000110111100100011 ;
        1887:  q   <=  32'b00111110001010001000001000101011 ;
        1888:  q   <=  32'b00111110001010001001010100110010 ;
        1889:  q   <=  32'b00111110001010001010100000111000 ;
        1890:  q   <=  32'b00111110001010001011101100111101 ;
        1891:  q   <=  32'b00111110001010001100111001000001 ;
        1892:  q   <=  32'b00111110001010001110000101000101 ;
        1893:  q   <=  32'b00111110001010001111010001001000 ;
        1894:  q   <=  32'b00111110001010010000011101001010 ;
        1895:  q   <=  32'b00111110001010010001101001001011 ;
        1896:  q   <=  32'b00111110001010010010110101001100 ;
        1897:  q   <=  32'b00111110001010010100000001001011 ;
        1898:  q   <=  32'b00111110001010010101001101001010 ;
        1899:  q   <=  32'b00111110001010010110011001001000 ;
        1900:  q   <=  32'b00111110001010010111100101000101 ;
        1901:  q   <=  32'b00111110001010011000110001000001 ;
        1902:  q   <=  32'b00111110001010011001111100111101 ;
        1903:  q   <=  32'b00111110001010011011001000111000 ;
        1904:  q   <=  32'b00111110001010011100010100110001 ;
        1905:  q   <=  32'b00111110001010011101100000101011 ;
        1906:  q   <=  32'b00111110001010011110101100100011 ;
        1907:  q   <=  32'b00111110001010011111111000011010 ;
        1908:  q   <=  32'b00111110001010100001000100010001 ;
        1909:  q   <=  32'b00111110001010100010010000000111 ;
        1910:  q   <=  32'b00111110001010100011011011111100 ;
        1911:  q   <=  32'b00111110001010100100100111110000 ;
        1912:  q   <=  32'b00111110001010100101110011100100 ;
        1913:  q   <=  32'b00111110001010100110111111010110 ;
        1914:  q   <=  32'b00111110001010101000001011001000 ;
        1915:  q   <=  32'b00111110001010101001010110111001 ;
        1916:  q   <=  32'b00111110001010101010100010101001 ;
        1917:  q   <=  32'b00111110001010101011101110011001 ;
        1918:  q   <=  32'b00111110001010101100111010000111 ;
        1919:  q   <=  32'b00111110001010101110000101110101 ;
        1920:  q   <=  32'b00111110001010101111010001100010 ;
        1921:  q   <=  32'b00111110001010110000011101001110 ;
        1922:  q   <=  32'b00111110001010110001101000111010 ;
        1923:  q   <=  32'b00111110001010110010110100100100 ;
        1924:  q   <=  32'b00111110001010110100000000001110 ;
        1925:  q   <=  32'b00111110001010110101001011110111 ;
        1926:  q   <=  32'b00111110001010110110010111011111 ;
        1927:  q   <=  32'b00111110001010110111100011000110 ;
        1928:  q   <=  32'b00111110001010111000101110101101 ;
        1929:  q   <=  32'b00111110001010111001111010010011 ;
        1930:  q   <=  32'b00111110001010111011000101111000 ;
        1931:  q   <=  32'b00111110001010111100010001011100 ;
        1932:  q   <=  32'b00111110001010111101011100111111 ;
        1933:  q   <=  32'b00111110001010111110101000100010 ;
        1934:  q   <=  32'b00111110001010111111110100000011 ;
        1935:  q   <=  32'b00111110001011000000111111100100 ;
        1936:  q   <=  32'b00111110001011000010001011000100 ;
        1937:  q   <=  32'b00111110001011000011010110100100 ;
        1938:  q   <=  32'b00111110001011000100100010000010 ;
        1939:  q   <=  32'b00111110001011000101101101100000 ;
        1940:  q   <=  32'b00111110001011000110111000111101 ;
        1941:  q   <=  32'b00111110001011001000000100011001 ;
        1942:  q   <=  32'b00111110001011001001001111110100 ;
        1943:  q   <=  32'b00111110001011001010011011001111 ;
        1944:  q   <=  32'b00111110001011001011100110101001 ;
        1945:  q   <=  32'b00111110001011001100110010000010 ;
        1946:  q   <=  32'b00111110001011001101111101011010 ;
        1947:  q   <=  32'b00111110001011001111001000110001 ;
        1948:  q   <=  32'b00111110001011010000010100001000 ;
        1949:  q   <=  32'b00111110001011010001011111011101 ;
        1950:  q   <=  32'b00111110001011010010101010110010 ;
        1951:  q   <=  32'b00111110001011010011110110000110 ;
        1952:  q   <=  32'b00111110001011010101000001011010 ;
        1953:  q   <=  32'b00111110001011010110001100101100 ;
        1954:  q   <=  32'b00111110001011010111010111111110 ;
        1955:  q   <=  32'b00111110001011011000100011001111 ;
        1956:  q   <=  32'b00111110001011011001101110011111 ;
        1957:  q   <=  32'b00111110001011011010111001101111 ;
        1958:  q   <=  32'b00111110001011011100000100111101 ;
        1959:  q   <=  32'b00111110001011011101010000001011 ;
        1960:  q   <=  32'b00111110001011011110011011011000 ;
        1961:  q   <=  32'b00111110001011011111100110100100 ;
        1962:  q   <=  32'b00111110001011100000110001110000 ;
        1963:  q   <=  32'b00111110001011100001111100111010 ;
        1964:  q   <=  32'b00111110001011100011001000000100 ;
        1965:  q   <=  32'b00111110001011100100010011001101 ;
        1966:  q   <=  32'b00111110001011100101011110010101 ;
        1967:  q   <=  32'b00111110001011100110101001011101 ;
        1968:  q   <=  32'b00111110001011100111110100100011 ;
        1969:  q   <=  32'b00111110001011101000111111101001 ;
        1970:  q   <=  32'b00111110001011101010001010101110 ;
        1971:  q   <=  32'b00111110001011101011010101110010 ;
        1972:  q   <=  32'b00111110001011101100100000110110 ;
        1973:  q   <=  32'b00111110001011101101101011111001 ;
        1974:  q   <=  32'b00111110001011101110110110111010 ;
        1975:  q   <=  32'b00111110001011110000000001111011 ;
        1976:  q   <=  32'b00111110001011110001001100111100 ;
        1977:  q   <=  32'b00111110001011110010010111111011 ;
        1978:  q   <=  32'b00111110001011110011100010111010 ;
        1979:  q   <=  32'b00111110001011110100101101111000 ;
        1980:  q   <=  32'b00111110001011110101111000110101 ;
        1981:  q   <=  32'b00111110001011110111000011110001 ;
        1982:  q   <=  32'b00111110001011111000001110101101 ;
        1983:  q   <=  32'b00111110001011111001011001101000 ;
        1984:  q   <=  32'b00111110001011111010100100100010 ;
        1985:  q   <=  32'b00111110001011111011101111011011 ;
        1986:  q   <=  32'b00111110001011111100111010010011 ;
        1987:  q   <=  32'b00111110001011111110000101001011 ;
        1988:  q   <=  32'b00111110001011111111010000000010 ;
        1989:  q   <=  32'b00111110001100000000011010111000 ;
        1990:  q   <=  32'b00111110001100000001100101101101 ;
        1991:  q   <=  32'b00111110001100000010110000100010 ;
        1992:  q   <=  32'b00111110001100000011111011010101 ;
        1993:  q   <=  32'b00111110001100000101000110001000 ;
        1994:  q   <=  32'b00111110001100000110010000111010 ;
        1995:  q   <=  32'b00111110001100000111011011101100 ;
        1996:  q   <=  32'b00111110001100001000100110011100 ;
        1997:  q   <=  32'b00111110001100001001110001001100 ;
        1998:  q   <=  32'b00111110001100001010111011111011 ;
        1999:  q   <=  32'b00111110001100001100000110101001 ;
        2000:  q   <=  32'b00111110001100001101010001010110 ;
        2001:  q   <=  32'b00111110001100001110011100000011 ;
        2002:  q   <=  32'b00111110001100001111100110101111 ;
        2003:  q   <=  32'b00111110001100010000110001011010 ;
        2004:  q   <=  32'b00111110001100010001111100000100 ;
        2005:  q   <=  32'b00111110001100010011000110101110 ;
        2006:  q   <=  32'b00111110001100010100010001010110 ;
        2007:  q   <=  32'b00111110001100010101011011111110 ;
        2008:  q   <=  32'b00111110001100010110100110100101 ;
        2009:  q   <=  32'b00111110001100010111110001001100 ;
        2010:  q   <=  32'b00111110001100011000111011110001 ;
        2011:  q   <=  32'b00111110001100011010000110010110 ;
        2012:  q   <=  32'b00111110001100011011010000111010 ;
        2013:  q   <=  32'b00111110001100011100011011011101 ;
        2014:  q   <=  32'b00111110001100011101100110000000 ;
        2015:  q   <=  32'b00111110001100011110110000100001 ;
        2016:  q   <=  32'b00111110001100011111111011000010 ;
        2017:  q   <=  32'b00111110001100100001000101100010 ;
        2018:  q   <=  32'b00111110001100100010010000000010 ;
        2019:  q   <=  32'b00111110001100100011011010100000 ;
        2020:  q   <=  32'b00111110001100100100100100111110 ;
        2021:  q   <=  32'b00111110001100100101101111011011 ;
        2022:  q   <=  32'b00111110001100100110111001110111 ;
        2023:  q   <=  32'b00111110001100101000000100010011 ;
        2024:  q   <=  32'b00111110001100101001001110101101 ;
        2025:  q   <=  32'b00111110001100101010011001000111 ;
        2026:  q   <=  32'b00111110001100101011100011100000 ;
        2027:  q   <=  32'b00111110001100101100101101111000 ;
        2028:  q   <=  32'b00111110001100101101111000010000 ;
        2029:  q   <=  32'b00111110001100101111000010100111 ;
        2030:  q   <=  32'b00111110001100110000001100111101 ;
        2031:  q   <=  32'b00111110001100110001010111010010 ;
        2032:  q   <=  32'b00111110001100110010100001100110 ;
        2033:  q   <=  32'b00111110001100110011101011111010 ;
        2034:  q   <=  32'b00111110001100110100110110001101 ;
        2035:  q   <=  32'b00111110001100110110000000011111 ;
        2036:  q   <=  32'b00111110001100110111001010110000 ;
        2037:  q   <=  32'b00111110001100111000010101000001 ;
        2038:  q   <=  32'b00111110001100111001011111010001 ;
        2039:  q   <=  32'b00111110001100111010101001100000 ;
        2040:  q   <=  32'b00111110001100111011110011101110 ;
        2041:  q   <=  32'b00111110001100111100111101111011 ;
        2042:  q   <=  32'b00111110001100111110001000001000 ;
        2043:  q   <=  32'b00111110001100111111010010010100 ;
        2044:  q   <=  32'b00111110001101000000011100011111 ;
        2045:  q   <=  32'b00111110001101000001100110101001 ;
        2046:  q   <=  32'b00111110001101000010110000110011 ;
        2047:  q   <=  32'b00111110001101000011111010111100 ;
        2048:  q   <=  32'b00111110001101000101000101000100 ;
        2049:  q   <=  32'b00111110001101000110001111001011 ;
        2050:  q   <=  32'b00111110001101000111011001010010 ;
        2051:  q   <=  32'b00111110001101001000100011010111 ;
        2052:  q   <=  32'b00111110001101001001101101011100 ;
        2053:  q   <=  32'b00111110001101001010110111100000 ;
        2054:  q   <=  32'b00111110001101001100000001100100 ;
        2055:  q   <=  32'b00111110001101001101001011100111 ;
        2056:  q   <=  32'b00111110001101001110010101101000 ;
        2057:  q   <=  32'b00111110001101001111011111101010 ;
        2058:  q   <=  32'b00111110001101010000101001101010 ;
        2059:  q   <=  32'b00111110001101010001110011101001 ;
        2060:  q   <=  32'b00111110001101010010111101101000 ;
        2061:  q   <=  32'b00111110001101010100000111100110 ;
        2062:  q   <=  32'b00111110001101010101010001100011 ;
        2063:  q   <=  32'b00111110001101010110011011100000 ;
        2064:  q   <=  32'b00111110001101010111100101011100 ;
        2065:  q   <=  32'b00111110001101011000101111010111 ;
        2066:  q   <=  32'b00111110001101011001111001010001 ;
        2067:  q   <=  32'b00111110001101011011000011001010 ;
        2068:  q   <=  32'b00111110001101011100001101000011 ;
        2069:  q   <=  32'b00111110001101011101010110111011 ;
        2070:  q   <=  32'b00111110001101011110100000110010 ;
        2071:  q   <=  32'b00111110001101011111101010101000 ;
        2072:  q   <=  32'b00111110001101100000110100011110 ;
        2073:  q   <=  32'b00111110001101100001111110010011 ;
        2074:  q   <=  32'b00111110001101100011001000000111 ;
        2075:  q   <=  32'b00111110001101100100010001111010 ;
        2076:  q   <=  32'b00111110001101100101011011101100 ;
        2077:  q   <=  32'b00111110001101100110100101011110 ;
        2078:  q   <=  32'b00111110001101100111101111001111 ;
        2079:  q   <=  32'b00111110001101101000111000111111 ;
        2080:  q   <=  32'b00111110001101101010000010101111 ;
        2081:  q   <=  32'b00111110001101101011001100011110 ;
        2082:  q   <=  32'b00111110001101101100010110001011 ;
        2083:  q   <=  32'b00111110001101101101011111111001 ;
        2084:  q   <=  32'b00111110001101101110101001100101 ;
        2085:  q   <=  32'b00111110001101101111110011010001 ;
        2086:  q   <=  32'b00111110001101110000111100111100 ;
        2087:  q   <=  32'b00111110001101110010000110100110 ;
        2088:  q   <=  32'b00111110001101110011010000001111 ;
        2089:  q   <=  32'b00111110001101110100011001111000 ;
        2090:  q   <=  32'b00111110001101110101100011011111 ;
        2091:  q   <=  32'b00111110001101110110101101000110 ;
        2092:  q   <=  32'b00111110001101110111110110101101 ;
        2093:  q   <=  32'b00111110001101111001000000010010 ;
        2094:  q   <=  32'b00111110001101111010001001110111 ;
        2095:  q   <=  32'b00111110001101111011010011011011 ;
        2096:  q   <=  32'b00111110001101111100011100111110 ;
        2097:  q   <=  32'b00111110001101111101100110100001 ;
        2098:  q   <=  32'b00111110001101111110110000000011 ;
        2099:  q   <=  32'b00111110001101111111111001100100 ;
        2100:  q   <=  32'b00111110001110000001000011000100 ;
        2101:  q   <=  32'b00111110001110000010001100100011 ;
        2102:  q   <=  32'b00111110001110000011010110000010 ;
        2103:  q   <=  32'b00111110001110000100011111100000 ;
        2104:  q   <=  32'b00111110001110000101101000111101 ;
        2105:  q   <=  32'b00111110001110000110110010011010 ;
        2106:  q   <=  32'b00111110001110000111111011110101 ;
        2107:  q   <=  32'b00111110001110001001000101010000 ;
        2108:  q   <=  32'b00111110001110001010001110101010 ;
        2109:  q   <=  32'b00111110001110001011011000000100 ;
        2110:  q   <=  32'b00111110001110001100100001011100 ;
        2111:  q   <=  32'b00111110001110001101101010110100 ;
        2112:  q   <=  32'b00111110001110001110110100001011 ;
        2113:  q   <=  32'b00111110001110001111111101100010 ;
        2114:  q   <=  32'b00111110001110010001000110110111 ;
        2115:  q   <=  32'b00111110001110010010010000001100 ;
        2116:  q   <=  32'b00111110001110010011011001100000 ;
        2117:  q   <=  32'b00111110001110010100100010110100 ;
        2118:  q   <=  32'b00111110001110010101101100000110 ;
        2119:  q   <=  32'b00111110001110010110110101011000 ;
        2120:  q   <=  32'b00111110001110010111111110101001 ;
        2121:  q   <=  32'b00111110001110011001000111111010 ;
        2122:  q   <=  32'b00111110001110011010010001001001 ;
        2123:  q   <=  32'b00111110001110011011011010011000 ;
        2124:  q   <=  32'b00111110001110011100100011100110 ;
        2125:  q   <=  32'b00111110001110011101101100110011 ;
        2126:  q   <=  32'b00111110001110011110110110000000 ;
        2127:  q   <=  32'b00111110001110011111111111001100 ;
        2128:  q   <=  32'b00111110001110100001001000010111 ;
        2129:  q   <=  32'b00111110001110100010010001100001 ;
        2130:  q   <=  32'b00111110001110100011011010101011 ;
        2131:  q   <=  32'b00111110001110100100100011110011 ;
        2132:  q   <=  32'b00111110001110100101101100111011 ;
        2133:  q   <=  32'b00111110001110100110110110000011 ;
        2134:  q   <=  32'b00111110001110100111111111001001 ;
        2135:  q   <=  32'b00111110001110101001001000001111 ;
        2136:  q   <=  32'b00111110001110101010010001010100 ;
        2137:  q   <=  32'b00111110001110101011011010011000 ;
        2138:  q   <=  32'b00111110001110101100100011011100 ;
        2139:  q   <=  32'b00111110001110101101101100011111 ;
        2140:  q   <=  32'b00111110001110101110110101100001 ;
        2141:  q   <=  32'b00111110001110101111111110100010 ;
        2142:  q   <=  32'b00111110001110110001000111100011 ;
        2143:  q   <=  32'b00111110001110110010010000100010 ;
        2144:  q   <=  32'b00111110001110110011011001100010 ;
        2145:  q   <=  32'b00111110001110110100100010100000 ;
        2146:  q   <=  32'b00111110001110110101101011011101 ;
        2147:  q   <=  32'b00111110001110110110110100011010 ;
        2148:  q   <=  32'b00111110001110110111111101010110 ;
        2149:  q   <=  32'b00111110001110111001000110010010 ;
        2150:  q   <=  32'b00111110001110111010001111001100 ;
        2151:  q   <=  32'b00111110001110111011011000000110 ;
        2152:  q   <=  32'b00111110001110111100100000111111 ;
        2153:  q   <=  32'b00111110001110111101101001110111 ;
        2154:  q   <=  32'b00111110001110111110110010101111 ;
        2155:  q   <=  32'b00111110001110111111111011100110 ;
        2156:  q   <=  32'b00111110001111000001000100011100 ;
        2157:  q   <=  32'b00111110001111000010001101010001 ;
        2158:  q   <=  32'b00111110001111000011010110000110 ;
        2159:  q   <=  32'b00111110001111000100011110111010 ;
        2160:  q   <=  32'b00111110001111000101100111101101 ;
        2161:  q   <=  32'b00111110001111000110110000011111 ;
        2162:  q   <=  32'b00111110001111000111111001010001 ;
        2163:  q   <=  32'b00111110001111001001000010000010 ;
        2164:  q   <=  32'b00111110001111001010001010110010 ;
        2165:  q   <=  32'b00111110001111001011010011100001 ;
        2166:  q   <=  32'b00111110001111001100011100010000 ;
        2167:  q   <=  32'b00111110001111001101100100111110 ;
        2168:  q   <=  32'b00111110001111001110101101101011 ;
        2169:  q   <=  32'b00111110001111001111110110010111 ;
        2170:  q   <=  32'b00111110001111010000111111000011 ;
        2171:  q   <=  32'b00111110001111010010000111101110 ;
        2172:  q   <=  32'b00111110001111010011010000011000 ;
        2173:  q   <=  32'b00111110001111010100011001000001 ;
        2174:  q   <=  32'b00111110001111010101100001101010 ;
        2175:  q   <=  32'b00111110001111010110101010010010 ;
        2176:  q   <=  32'b00111110001111010111110010111001 ;
        2177:  q   <=  32'b00111110001111011000111011100000 ;
        2178:  q   <=  32'b00111110001111011010000100000101 ;
        2179:  q   <=  32'b00111110001111011011001100101010 ;
        2180:  q   <=  32'b00111110001111011100010101001111 ;
        2181:  q   <=  32'b00111110001111011101011101110010 ;
        2182:  q   <=  32'b00111110001111011110100110010101 ;
        2183:  q   <=  32'b00111110001111011111101110110111 ;
        2184:  q   <=  32'b00111110001111100000110111011000 ;
        2185:  q   <=  32'b00111110001111100001111111111001 ;
        2186:  q   <=  32'b00111110001111100011001000011001 ;
        2187:  q   <=  32'b00111110001111100100010000111000 ;
        2188:  q   <=  32'b00111110001111100101011001010110 ;
        2189:  q   <=  32'b00111110001111100110100001110100 ;
        2190:  q   <=  32'b00111110001111100111101010010000 ;
        2191:  q   <=  32'b00111110001111101000110010101101 ;
        2192:  q   <=  32'b00111110001111101001111011001000 ;
        2193:  q   <=  32'b00111110001111101011000011100011 ;
        2194:  q   <=  32'b00111110001111101100001011111101 ;
        2195:  q   <=  32'b00111110001111101101010100010110 ;
        2196:  q   <=  32'b00111110001111101110011100101110 ;
        2197:  q   <=  32'b00111110001111101111100101000110 ;
        2198:  q   <=  32'b00111110001111110000101101011101 ;
        2199:  q   <=  32'b00111110001111110001110101110011 ;
        2200:  q   <=  32'b00111110001111110010111110001001 ;
        2201:  q   <=  32'b00111110001111110100000110011101 ;
        2202:  q   <=  32'b00111110001111110101001110110001 ;
        2203:  q   <=  32'b00111110001111110110010111000101 ;
        2204:  q   <=  32'b00111110001111110111011111010111 ;
        2205:  q   <=  32'b00111110001111111000100111101001 ;
        2206:  q   <=  32'b00111110001111111001101111111010 ;
        2207:  q   <=  32'b00111110001111111010111000001011 ;
        2208:  q   <=  32'b00111110001111111100000000011010 ;
        2209:  q   <=  32'b00111110001111111101001000101001 ;
        2210:  q   <=  32'b00111110001111111110010000110111 ;
        2211:  q   <=  32'b00111110001111111111011001000101 ;
        2212:  q   <=  32'b00111110010000000000100001010001 ;
        2213:  q   <=  32'b00111110010000000001101001011101 ;
        2214:  q   <=  32'b00111110010000000010110001101000 ;
        2215:  q   <=  32'b00111110010000000011111001110011 ;
        2216:  q   <=  32'b00111110010000000101000001111101 ;
        2217:  q   <=  32'b00111110010000000110001010000110 ;
        2218:  q   <=  32'b00111110010000000111010010001110 ;
        2219:  q   <=  32'b00111110010000001000011010010110 ;
        2220:  q   <=  32'b00111110010000001001100010011100 ;
        2221:  q   <=  32'b00111110010000001010101010100011 ;
        2222:  q   <=  32'b00111110010000001011110010101000 ;
        2223:  q   <=  32'b00111110010000001100111010101101 ;
        2224:  q   <=  32'b00111110010000001110000010110001 ;
        2225:  q   <=  32'b00111110010000001111001010110100 ;
        2226:  q   <=  32'b00111110010000010000010010110110 ;
        2227:  q   <=  32'b00111110010000010001011010111000 ;
        2228:  q   <=  32'b00111110010000010010100010111001 ;
        2229:  q   <=  32'b00111110010000010011101010111001 ;
        2230:  q   <=  32'b00111110010000010100110010111001 ;
        2231:  q   <=  32'b00111110010000010101111010111000 ;
        2232:  q   <=  32'b00111110010000010111000010110110 ;
        2233:  q   <=  32'b00111110010000011000001010110011 ;
        2234:  q   <=  32'b00111110010000011001010010110000 ;
        2235:  q   <=  32'b00111110010000011010011010101100 ;
        2236:  q   <=  32'b00111110010000011011100010100111 ;
        2237:  q   <=  32'b00111110010000011100101010100001 ;
        2238:  q   <=  32'b00111110010000011101110010011011 ;
        2239:  q   <=  32'b00111110010000011110111010010100 ;
        2240:  q   <=  32'b00111110010000100000000010001100 ;
        2241:  q   <=  32'b00111110010000100001001010000100 ;
        2242:  q   <=  32'b00111110010000100010010001111010 ;
        2243:  q   <=  32'b00111110010000100011011001110001 ;
        2244:  q   <=  32'b00111110010000100100100001100110 ;
        2245:  q   <=  32'b00111110010000100101101001011011 ;
        2246:  q   <=  32'b00111110010000100110110001001111 ;
        2247:  q   <=  32'b00111110010000100111111001000010 ;
        2248:  q   <=  32'b00111110010000101001000000110100 ;
        2249:  q   <=  32'b00111110010000101010001000100110 ;
        2250:  q   <=  32'b00111110010000101011010000010111 ;
        2251:  q   <=  32'b00111110010000101100011000000111 ;
        2252:  q   <=  32'b00111110010000101101011111110111 ;
        2253:  q   <=  32'b00111110010000101110100111100110 ;
        2254:  q   <=  32'b00111110010000101111101111010100 ;
        2255:  q   <=  32'b00111110010000110000110111000001 ;
        2256:  q   <=  32'b00111110010000110001111110101110 ;
        2257:  q   <=  32'b00111110010000110011000110011010 ;
        2258:  q   <=  32'b00111110010000110100001110000101 ;
        2259:  q   <=  32'b00111110010000110101010101110000 ;
        2260:  q   <=  32'b00111110010000110110011101011001 ;
        2261:  q   <=  32'b00111110010000110111100101000010 ;
        2262:  q   <=  32'b00111110010000111000101100101011 ;
        2263:  q   <=  32'b00111110010000111001110100010010 ;
        2264:  q   <=  32'b00111110010000111010111011111001 ;
        2265:  q   <=  32'b00111110010000111100000011100000 ;
        2266:  q   <=  32'b00111110010000111101001011000101 ;
        2267:  q   <=  32'b00111110010000111110010010101010 ;
        2268:  q   <=  32'b00111110010000111111011010001110 ;
        2269:  q   <=  32'b00111110010001000000100001110001 ;
        2270:  q   <=  32'b00111110010001000001101001010100 ;
        2271:  q   <=  32'b00111110010001000010110000110110 ;
        2272:  q   <=  32'b00111110010001000011111000010111 ;
        2273:  q   <=  32'b00111110010001000100111111110111 ;
        2274:  q   <=  32'b00111110010001000110000111010111 ;
        2275:  q   <=  32'b00111110010001000111001110110110 ;
        2276:  q   <=  32'b00111110010001001000010110010100 ;
        2277:  q   <=  32'b00111110010001001001011101110010 ;
        2278:  q   <=  32'b00111110010001001010100101001111 ;
        2279:  q   <=  32'b00111110010001001011101100101011 ;
        2280:  q   <=  32'b00111110010001001100110100000110 ;
        2281:  q   <=  32'b00111110010001001101111011100001 ;
        2282:  q   <=  32'b00111110010001001111000010111011 ;
        2283:  q   <=  32'b00111110010001010000001010010100 ;
        2284:  q   <=  32'b00111110010001010001010001101101 ;
        2285:  q   <=  32'b00111110010001010010011001000100 ;
        2286:  q   <=  32'b00111110010001010011100000011011 ;
        2287:  q   <=  32'b00111110010001010100100111110010 ;
        2288:  q   <=  32'b00111110010001010101101111001000 ;
        2289:  q   <=  32'b00111110010001010110110110011100 ;
        2290:  q   <=  32'b00111110010001010111111101110001 ;
        2291:  q   <=  32'b00111110010001011001000101000100 ;
        2292:  q   <=  32'b00111110010001011010001100010111 ;
        2293:  q   <=  32'b00111110010001011011010011101001 ;
        2294:  q   <=  32'b00111110010001011100011010111011 ;
        2295:  q   <=  32'b00111110010001011101100010001011 ;
        2296:  q   <=  32'b00111110010001011110101001011011 ;
        2297:  q   <=  32'b00111110010001011111110000101010 ;
        2298:  q   <=  32'b00111110010001100000110111111001 ;
        2299:  q   <=  32'b00111110010001100001111111000111 ;
        2300:  q   <=  32'b00111110010001100011000110010100 ;
        2301:  q   <=  32'b00111110010001100100001101100000 ;
        2302:  q   <=  32'b00111110010001100101010100101100 ;
        2303:  q   <=  32'b00111110010001100110011011110111 ;
        2304:  q   <=  32'b00111110010001100111100011000001 ;
        2305:  q   <=  32'b00111110010001101000101010001011 ;
        2306:  q   <=  32'b00111110010001101001110001010100 ;
        2307:  q   <=  32'b00111110010001101010111000011100 ;
        2308:  q   <=  32'b00111110010001101011111111100011 ;
        2309:  q   <=  32'b00111110010001101101000110101010 ;
        2310:  q   <=  32'b00111110010001101110001101110000 ;
        2311:  q   <=  32'b00111110010001101111010100110101 ;
        2312:  q   <=  32'b00111110010001110000011011111010 ;
        2313:  q   <=  32'b00111110010001110001100010111110 ;
        2314:  q   <=  32'b00111110010001110010101010000001 ;
        2315:  q   <=  32'b00111110010001110011110001000011 ;
        2316:  q   <=  32'b00111110010001110100111000000101 ;
        2317:  q   <=  32'b00111110010001110101111111000110 ;
        2318:  q   <=  32'b00111110010001110111000110000110 ;
        2319:  q   <=  32'b00111110010001111000001101000110 ;
        2320:  q   <=  32'b00111110010001111001010100000101 ;
        2321:  q   <=  32'b00111110010001111010011011000011 ;
        2322:  q   <=  32'b00111110010001111011100010000001 ;
        2323:  q   <=  32'b00111110010001111100101000111101 ;
        2324:  q   <=  32'b00111110010001111101101111111001 ;
        2325:  q   <=  32'b00111110010001111110110110110101 ;
        2326:  q   <=  32'b00111110010001111111111101101111 ;
        2327:  q   <=  32'b00111110010010000001000100101001 ;
        2328:  q   <=  32'b00111110010010000010001011100011 ;
        2329:  q   <=  32'b00111110010010000011010010011011 ;
        2330:  q   <=  32'b00111110010010000100011001010011 ;
        2331:  q   <=  32'b00111110010010000101100000001010 ;
        2332:  q   <=  32'b00111110010010000110100111000001 ;
        2333:  q   <=  32'b00111110010010000111101101110110 ;
        2334:  q   <=  32'b00111110010010001000110100101011 ;
        2335:  q   <=  32'b00111110010010001001111011100000 ;
        2336:  q   <=  32'b00111110010010001011000010010011 ;
        2337:  q   <=  32'b00111110010010001100001001000110 ;
        2338:  q   <=  32'b00111110010010001101001111111000 ;
        2339:  q   <=  32'b00111110010010001110010110101010 ;
        2340:  q   <=  32'b00111110010010001111011101011011 ;
        2341:  q   <=  32'b00111110010010010000100100001011 ;
        2342:  q   <=  32'b00111110010010010001101010111010 ;
        2343:  q   <=  32'b00111110010010010010110001101001 ;
        2344:  q   <=  32'b00111110010010010011111000010111 ;
        2345:  q   <=  32'b00111110010010010100111111000100 ;
        2346:  q   <=  32'b00111110010010010110000101110001 ;
        2347:  q   <=  32'b00111110010010010111001100011100 ;
        2348:  q   <=  32'b00111110010010011000010011001000 ;
        2349:  q   <=  32'b00111110010010011001011001110010 ;
        2350:  q   <=  32'b00111110010010011010100000011100 ;
        2351:  q   <=  32'b00111110010010011011100111000101 ;
        2352:  q   <=  32'b00111110010010011100101101101101 ;
        2353:  q   <=  32'b00111110010010011101110100010101 ;
        2354:  q   <=  32'b00111110010010011110111010111100 ;
        2355:  q   <=  32'b00111110010010100000000001100010 ;
        2356:  q   <=  32'b00111110010010100001001000001000 ;
        2357:  q   <=  32'b00111110010010100010001110101100 ;
        2358:  q   <=  32'b00111110010010100011010101010001 ;
        2359:  q   <=  32'b00111110010010100100011011110100 ;
        2360:  q   <=  32'b00111110010010100101100010010111 ;
        2361:  q   <=  32'b00111110010010100110101000111001 ;
        2362:  q   <=  32'b00111110010010100111101111011010 ;
        2363:  q   <=  32'b00111110010010101000110101111011 ;
        2364:  q   <=  32'b00111110010010101001111100011011 ;
        2365:  q   <=  32'b00111110010010101011000010111010 ;
        2366:  q   <=  32'b00111110010010101100001001011001 ;
        2367:  q   <=  32'b00111110010010101101001111110111 ;
        2368:  q   <=  32'b00111110010010101110010110010100 ;
        2369:  q   <=  32'b00111110010010101111011100110000 ;
        2370:  q   <=  32'b00111110010010110000100011001100 ;
        2371:  q   <=  32'b00111110010010110001101001100111 ;
        2372:  q   <=  32'b00111110010010110010110000000001 ;
        2373:  q   <=  32'b00111110010010110011110110011011 ;
        2374:  q   <=  32'b00111110010010110100111100110100 ;
        2375:  q   <=  32'b00111110010010110110000011001100 ;
        2376:  q   <=  32'b00111110010010110111001001100100 ;
        2377:  q   <=  32'b00111110010010111000001111111011 ;
        2378:  q   <=  32'b00111110010010111001010110010001 ;
        2379:  q   <=  32'b00111110010010111010011100100111 ;
        2380:  q   <=  32'b00111110010010111011100010111011 ;
        2381:  q   <=  32'b00111110010010111100101001010000 ;
        2382:  q   <=  32'b00111110010010111101101111100011 ;
        2383:  q   <=  32'b00111110010010111110110101110110 ;
        2384:  q   <=  32'b00111110010010111111111100001000 ;
        2385:  q   <=  32'b00111110010011000001000010011001 ;
        2386:  q   <=  32'b00111110010011000010001000101010 ;
        2387:  q   <=  32'b00111110010011000011001110111010 ;
        2388:  q   <=  32'b00111110010011000100010101001001 ;
        2389:  q   <=  32'b00111110010011000101011011010111 ;
        2390:  q   <=  32'b00111110010011000110100001100101 ;
        2391:  q   <=  32'b00111110010011000111100111110011 ;
        2392:  q   <=  32'b00111110010011001000101101111111 ;
        2393:  q   <=  32'b00111110010011001001110100001011 ;
        2394:  q   <=  32'b00111110010011001010111010010110 ;
        2395:  q   <=  32'b00111110010011001100000000100000 ;
        2396:  q   <=  32'b00111110010011001101000110101010 ;
        2397:  q   <=  32'b00111110010011001110001100110011 ;
        2398:  q   <=  32'b00111110010011001111010010111011 ;
        2399:  q   <=  32'b00111110010011010000011001000011 ;
        2400:  q   <=  32'b00111110010011010001011111001010 ;
        2401:  q   <=  32'b00111110010011010010100101010000 ;
        2402:  q   <=  32'b00111110010011010011101011010110 ;
        2403:  q   <=  32'b00111110010011010100110001011011 ;
        2404:  q   <=  32'b00111110010011010101110111011111 ;
        2405:  q   <=  32'b00111110010011010110111101100010 ;
        2406:  q   <=  32'b00111110010011011000000011100101 ;
        2407:  q   <=  32'b00111110010011011001001001100111 ;
        2408:  q   <=  32'b00111110010011011010001111101001 ;
        2409:  q   <=  32'b00111110010011011011010101101010 ;
        2410:  q   <=  32'b00111110010011011100011011101010 ;
        2411:  q   <=  32'b00111110010011011101100001101001 ;
        2412:  q   <=  32'b00111110010011011110100111101000 ;
        2413:  q   <=  32'b00111110010011011111101101100110 ;
        2414:  q   <=  32'b00111110010011100000110011100011 ;
        2415:  q   <=  32'b00111110010011100001111001100000 ;
        2416:  q   <=  32'b00111110010011100010111111011011 ;
        2417:  q   <=  32'b00111110010011100100000101010111 ;
        2418:  q   <=  32'b00111110010011100101001011010001 ;
        2419:  q   <=  32'b00111110010011100110010001001011 ;
        2420:  q   <=  32'b00111110010011100111010111000100 ;
        2421:  q   <=  32'b00111110010011101000011100111101 ;
        2422:  q   <=  32'b00111110010011101001100010110101 ;
        2423:  q   <=  32'b00111110010011101010101000101100 ;
        2424:  q   <=  32'b00111110010011101011101110100010 ;
        2425:  q   <=  32'b00111110010011101100110100011000 ;
        2426:  q   <=  32'b00111110010011101101111010001101 ;
        2427:  q   <=  32'b00111110010011101111000000000001 ;
        2428:  q   <=  32'b00111110010011110000000101110101 ;
        2429:  q   <=  32'b00111110010011110001001011101000 ;
        2430:  q   <=  32'b00111110010011110010010001011010 ;
        2431:  q   <=  32'b00111110010011110011010111001100 ;
        2432:  q   <=  32'b00111110010011110100011100111101 ;
        2433:  q   <=  32'b00111110010011110101100010101101 ;
        2434:  q   <=  32'b00111110010011110110101000011101 ;
        2435:  q   <=  32'b00111110010011110111101110001100 ;
        2436:  q   <=  32'b00111110010011111000110011111010 ;
        2437:  q   <=  32'b00111110010011111001111001101000 ;
        2438:  q   <=  32'b00111110010011111010111111010100 ;
        2439:  q   <=  32'b00111110010011111100000101000001 ;
        2440:  q   <=  32'b00111110010011111101001010101100 ;
        2441:  q   <=  32'b00111110010011111110010000010111 ;
        2442:  q   <=  32'b00111110010011111111010110000001 ;
        2443:  q   <=  32'b00111110010100000000011011101010 ;
        2444:  q   <=  32'b00111110010100000001100001010011 ;
        2445:  q   <=  32'b00111110010100000010100110111011 ;
        2446:  q   <=  32'b00111110010100000011101100100011 ;
        2447:  q   <=  32'b00111110010100000100110010001001 ;
        2448:  q   <=  32'b00111110010100000101110111101111 ;
        2449:  q   <=  32'b00111110010100000110111101010101 ;
        2450:  q   <=  32'b00111110010100001000000010111010 ;
        2451:  q   <=  32'b00111110010100001001001000011110 ;
        2452:  q   <=  32'b00111110010100001010001110000001 ;
        2453:  q   <=  32'b00111110010100001011010011100011 ;
        2454:  q   <=  32'b00111110010100001100011001000101 ;
        2455:  q   <=  32'b00111110010100001101011110100111 ;
        2456:  q   <=  32'b00111110010100001110100100000111 ;
        2457:  q   <=  32'b00111110010100001111101001100111 ;
        2458:  q   <=  32'b00111110010100010000101111000110 ;
        2459:  q   <=  32'b00111110010100010001110100100101 ;
        2460:  q   <=  32'b00111110010100010010111010000011 ;
        2461:  q   <=  32'b00111110010100010011111111100000 ;
        2462:  q   <=  32'b00111110010100010101000100111101 ;
        2463:  q   <=  32'b00111110010100010110001010011001 ;
        2464:  q   <=  32'b00111110010100010111001111110100 ;
        2465:  q   <=  32'b00111110010100011000010101001110 ;
        2466:  q   <=  32'b00111110010100011001011010101000 ;
        2467:  q   <=  32'b00111110010100011010100000000001 ;
        2468:  q   <=  32'b00111110010100011011100101011010 ;
        2469:  q   <=  32'b00111110010100011100101010110001 ;
        2470:  q   <=  32'b00111110010100011101110000001001 ;
        2471:  q   <=  32'b00111110010100011110110101011111 ;
        2472:  q   <=  32'b00111110010100011111111010110101 ;
        2473:  q   <=  32'b00111110010100100001000000001010 ;
        2474:  q   <=  32'b00111110010100100010000101011110 ;
        2475:  q   <=  32'b00111110010100100011001010110010 ;
        2476:  q   <=  32'b00111110010100100100010000000101 ;
        2477:  q   <=  32'b00111110010100100101010101010111 ;
        2478:  q   <=  32'b00111110010100100110011010101001 ;
        2479:  q   <=  32'b00111110010100100111011111111010 ;
        2480:  q   <=  32'b00111110010100101000100101001011 ;
        2481:  q   <=  32'b00111110010100101001101010011010 ;
        2482:  q   <=  32'b00111110010100101010101111101001 ;
        2483:  q   <=  32'b00111110010100101011110100111000 ;
        2484:  q   <=  32'b00111110010100101100111010000101 ;
        2485:  q   <=  32'b00111110010100101101111111010010 ;
        2486:  q   <=  32'b00111110010100101111000100011111 ;
        2487:  q   <=  32'b00111110010100110000001001101010 ;
        2488:  q   <=  32'b00111110010100110001001110110101 ;
        2489:  q   <=  32'b00111110010100110010010100000000 ;
        2490:  q   <=  32'b00111110010100110011011001001001 ;
        2491:  q   <=  32'b00111110010100110100011110010010 ;
        2492:  q   <=  32'b00111110010100110101100011011010 ;
        2493:  q   <=  32'b00111110010100110110101000100010 ;
        2494:  q   <=  32'b00111110010100110111101101101001 ;
        2495:  q   <=  32'b00111110010100111000110010101111 ;
        2496:  q   <=  32'b00111110010100111001110111110101 ;
        2497:  q   <=  32'b00111110010100111010111100111010 ;
        2498:  q   <=  32'b00111110010100111100000001111110 ;
        2499:  q   <=  32'b00111110010100111101000111000010 ;
        2500:  q   <=  32'b00111110010100111110001100000101 ;
        2501:  q   <=  32'b00111110010100111111010001000111 ;
        2502:  q   <=  32'b00111110010101000000010110001000 ;
        2503:  q   <=  32'b00111110010101000001011011001001 ;
        2504:  q   <=  32'b00111110010101000010100000001010 ;
        2505:  q   <=  32'b00111110010101000011100101001001 ;
        2506:  q   <=  32'b00111110010101000100101010001000 ;
        2507:  q   <=  32'b00111110010101000101101111000110 ;
        2508:  q   <=  32'b00111110010101000110110100000100 ;
        2509:  q   <=  32'b00111110010101000111111001000001 ;
        2510:  q   <=  32'b00111110010101001000111101111101 ;
        2511:  q   <=  32'b00111110010101001010000010111001 ;
        2512:  q   <=  32'b00111110010101001011000111110011 ;
        2513:  q   <=  32'b00111110010101001100001100101110 ;
        2514:  q   <=  32'b00111110010101001101010001100111 ;
        2515:  q   <=  32'b00111110010101001110010110100000 ;
        2516:  q   <=  32'b00111110010101001111011011011000 ;
        2517:  q   <=  32'b00111110010101010000100000010000 ;
        2518:  q   <=  32'b00111110010101010001100101000111 ;
        2519:  q   <=  32'b00111110010101010010101001111101 ;
        2520:  q   <=  32'b00111110010101010011101110110011 ;
        2521:  q   <=  32'b00111110010101010100110011101000 ;
        2522:  q   <=  32'b00111110010101010101111000011100 ;
        2523:  q   <=  32'b00111110010101010110111101001111 ;
        2524:  q   <=  32'b00111110010101011000000010000010 ;
        2525:  q   <=  32'b00111110010101011001000110110100 ;
        2526:  q   <=  32'b00111110010101011010001011100110 ;
        2527:  q   <=  32'b00111110010101011011010000010111 ;
        2528:  q   <=  32'b00111110010101011100010101000111 ;
        2529:  q   <=  32'b00111110010101011101011001110111 ;
        2530:  q   <=  32'b00111110010101011110011110100110 ;
        2531:  q   <=  32'b00111110010101011111100011010100 ;
        2532:  q   <=  32'b00111110010101100000101000000010 ;
        2533:  q   <=  32'b00111110010101100001101100101110 ;
        2534:  q   <=  32'b00111110010101100010110001011011 ;
        2535:  q   <=  32'b00111110010101100011110110000110 ;
        2536:  q   <=  32'b00111110010101100100111010110001 ;
        2537:  q   <=  32'b00111110010101100101111111011011 ;
        2538:  q   <=  32'b00111110010101100111000100000101 ;
        2539:  q   <=  32'b00111110010101101000001000101110 ;
        2540:  q   <=  32'b00111110010101101001001101010110 ;
        2541:  q   <=  32'b00111110010101101010010001111110 ;
        2542:  q   <=  32'b00111110010101101011010110100101 ;
        2543:  q   <=  32'b00111110010101101100011011001011 ;
        2544:  q   <=  32'b00111110010101101101011111110001 ;
        2545:  q   <=  32'b00111110010101101110100100010110 ;
        2546:  q   <=  32'b00111110010101101111101000111010 ;
        2547:  q   <=  32'b00111110010101110000101101011110 ;
        2548:  q   <=  32'b00111110010101110001110010000001 ;
        2549:  q   <=  32'b00111110010101110010110110100011 ;
        2550:  q   <=  32'b00111110010101110011111011000101 ;
        2551:  q   <=  32'b00111110010101110100111111100110 ;
        2552:  q   <=  32'b00111110010101110110000100000110 ;
        2553:  q   <=  32'b00111110010101110111001000100110 ;
        2554:  q   <=  32'b00111110010101111000001101000101 ;
        2555:  q   <=  32'b00111110010101111001010001100011 ;
        2556:  q   <=  32'b00111110010101111010010110000001 ;
        2557:  q   <=  32'b00111110010101111011011010011110 ;
        2558:  q   <=  32'b00111110010101111100011110111010 ;
        2559:  q   <=  32'b00111110010101111101100011010110 ;
        2560:  q   <=  32'b00111110010101111110100111110001 ;
        2561:  q   <=  32'b00111110010101111111101100001100 ;
        2562:  q   <=  32'b00111110010110000000110000100110 ;
        2563:  q   <=  32'b00111110010110000001110100111111 ;
        2564:  q   <=  32'b00111110010110000010111001010111 ;
        2565:  q   <=  32'b00111110010110000011111101101111 ;
        2566:  q   <=  32'b00111110010110000101000010000110 ;
        2567:  q   <=  32'b00111110010110000110000110011101 ;
        2568:  q   <=  32'b00111110010110000111001010110010 ;
        2569:  q   <=  32'b00111110010110001000001111001000 ;
        2570:  q   <=  32'b00111110010110001001010011011100 ;
        2571:  q   <=  32'b00111110010110001010010111110000 ;
        2572:  q   <=  32'b00111110010110001011011100000011 ;
        2573:  q   <=  32'b00111110010110001100100000010110 ;
        2574:  q   <=  32'b00111110010110001101100100101000 ;
        2575:  q   <=  32'b00111110010110001110101000111001 ;
        2576:  q   <=  32'b00111110010110001111101101001001 ;
        2577:  q   <=  32'b00111110010110010000110001011001 ;
        2578:  q   <=  32'b00111110010110010001110101101001 ;
        2579:  q   <=  32'b00111110010110010010111001110111 ;
        2580:  q   <=  32'b00111110010110010011111110000101 ;
        2581:  q   <=  32'b00111110010110010101000010010010 ;
        2582:  q   <=  32'b00111110010110010110000110011111 ;
        2583:  q   <=  32'b00111110010110010111001010101011 ;
        2584:  q   <=  32'b00111110010110011000001110110110 ;
        2585:  q   <=  32'b00111110010110011001010011000001 ;
        2586:  q   <=  32'b00111110010110011010010111001011 ;
        2587:  q   <=  32'b00111110010110011011011011010101 ;
        2588:  q   <=  32'b00111110010110011100011111011101 ;
        2589:  q   <=  32'b00111110010110011101100011100101 ;
        2590:  q   <=  32'b00111110010110011110100111101101 ;
        2591:  q   <=  32'b00111110010110011111101011110100 ;
        2592:  q   <=  32'b00111110010110100000101111111010 ;
        2593:  q   <=  32'b00111110010110100001110011111111 ;
        2594:  q   <=  32'b00111110010110100010111000000100 ;
        2595:  q   <=  32'b00111110010110100011111100001000 ;
        2596:  q   <=  32'b00111110010110100101000000001100 ;
        2597:  q   <=  32'b00111110010110100110000100001111 ;
        2598:  q   <=  32'b00111110010110100111001000010001 ;
        2599:  q   <=  32'b00111110010110101000001100010010 ;
        2600:  q   <=  32'b00111110010110101001010000010011 ;
        2601:  q   <=  32'b00111110010110101010010100010100 ;
        2602:  q   <=  32'b00111110010110101011011000010011 ;
        2603:  q   <=  32'b00111110010110101100011100010010 ;
        2604:  q   <=  32'b00111110010110101101100000010001 ;
        2605:  q   <=  32'b00111110010110101110100100001110 ;
        2606:  q   <=  32'b00111110010110101111101000001011 ;
        2607:  q   <=  32'b00111110010110110000101100001000 ;
        2608:  q   <=  32'b00111110010110110001110000000011 ;
        2609:  q   <=  32'b00111110010110110010110011111111 ;
        2610:  q   <=  32'b00111110010110110011110111111001 ;
        2611:  q   <=  32'b00111110010110110100111011110011 ;
        2612:  q   <=  32'b00111110010110110101111111101100 ;
        2613:  q   <=  32'b00111110010110110111000011100100 ;
        2614:  q   <=  32'b00111110010110111000000111011100 ;
        2615:  q   <=  32'b00111110010110111001001011010011 ;
        2616:  q   <=  32'b00111110010110111010001111001010 ;
        2617:  q   <=  32'b00111110010110111011010011000000 ;
        2618:  q   <=  32'b00111110010110111100010110110101 ;
        2619:  q   <=  32'b00111110010110111101011010101010 ;
        2620:  q   <=  32'b00111110010110111110011110011110 ;
        2621:  q   <=  32'b00111110010110111111100010010001 ;
        2622:  q   <=  32'b00111110010111000000100110000100 ;
        2623:  q   <=  32'b00111110010111000001101001110110 ;
        2624:  q   <=  32'b00111110010111000010101101100111 ;
        2625:  q   <=  32'b00111110010111000011110001011000 ;
        2626:  q   <=  32'b00111110010111000100110101001000 ;
        2627:  q   <=  32'b00111110010111000101111000110111 ;
        2628:  q   <=  32'b00111110010111000110111100100110 ;
        2629:  q   <=  32'b00111110010111001000000000010100 ;
        2630:  q   <=  32'b00111110010111001001000100000010 ;
        2631:  q   <=  32'b00111110010111001010000111101111 ;
        2632:  q   <=  32'b00111110010111001011001011011011 ;
        2633:  q   <=  32'b00111110010111001100001111000110 ;
        2634:  q   <=  32'b00111110010111001101010010110001 ;
        2635:  q   <=  32'b00111110010111001110010110011100 ;
        2636:  q   <=  32'b00111110010111001111011010000101 ;
        2637:  q   <=  32'b00111110010111010000011101101110 ;
        2638:  q   <=  32'b00111110010111010001100001010111 ;
        2639:  q   <=  32'b00111110010111010010100100111110 ;
        2640:  q   <=  32'b00111110010111010011101000100101 ;
        2641:  q   <=  32'b00111110010111010100101100001100 ;
        2642:  q   <=  32'b00111110010111010101101111110010 ;
        2643:  q   <=  32'b00111110010111010110110011010111 ;
        2644:  q   <=  32'b00111110010111010111110110111011 ;
        2645:  q   <=  32'b00111110010111011000111010011111 ;
        2646:  q   <=  32'b00111110010111011001111110000010 ;
        2647:  q   <=  32'b00111110010111011011000001100101 ;
        2648:  q   <=  32'b00111110010111011100000101000111 ;
        2649:  q   <=  32'b00111110010111011101001000101000 ;
        2650:  q   <=  32'b00111110010111011110001100001001 ;
        2651:  q   <=  32'b00111110010111011111001111101001 ;
        2652:  q   <=  32'b00111110010111100000010011001000 ;
        2653:  q   <=  32'b00111110010111100001010110100111 ;
        2654:  q   <=  32'b00111110010111100010011010000101 ;
        2655:  q   <=  32'b00111110010111100011011101100011 ;
        2656:  q   <=  32'b00111110010111100100100000111111 ;
        2657:  q   <=  32'b00111110010111100101100100011100 ;
        2658:  q   <=  32'b00111110010111100110100111110111 ;
        2659:  q   <=  32'b00111110010111100111101011010010 ;
        2660:  q   <=  32'b00111110010111101000101110101100 ;
        2661:  q   <=  32'b00111110010111101001110010000110 ;
        2662:  q   <=  32'b00111110010111101010110101011111 ;
        2663:  q   <=  32'b00111110010111101011111000110111 ;
        2664:  q   <=  32'b00111110010111101100111100001111 ;
        2665:  q   <=  32'b00111110010111101101111111100110 ;
        2666:  q   <=  32'b00111110010111101111000010111100 ;
        2667:  q   <=  32'b00111110010111110000000110010010 ;
        2668:  q   <=  32'b00111110010111110001001001100111 ;
        2669:  q   <=  32'b00111110010111110010001100111100 ;
        2670:  q   <=  32'b00111110010111110011010000010000 ;
        2671:  q   <=  32'b00111110010111110100010011100011 ;
        2672:  q   <=  32'b00111110010111110101010110110110 ;
        2673:  q   <=  32'b00111110010111110110011010001000 ;
        2674:  q   <=  32'b00111110010111110111011101011001 ;
        2675:  q   <=  32'b00111110010111111000100000101010 ;
        2676:  q   <=  32'b00111110010111111001100011111010 ;
        2677:  q   <=  32'b00111110010111111010100111001001 ;
        2678:  q   <=  32'b00111110010111111011101010011000 ;
        2679:  q   <=  32'b00111110010111111100101101100110 ;
        2680:  q   <=  32'b00111110010111111101110000110100 ;
        2681:  q   <=  32'b00111110010111111110110100000001 ;
        2682:  q   <=  32'b00111110010111111111110111001101 ;
        2683:  q   <=  32'b00111110011000000000111010011001 ;
        2684:  q   <=  32'b00111110011000000001111101100100 ;
        2685:  q   <=  32'b00111110011000000011000000101110 ;
        2686:  q   <=  32'b00111110011000000100000011111000 ;
        2687:  q   <=  32'b00111110011000000101000111000001 ;
        2688:  q   <=  32'b00111110011000000110001010001001 ;
        2689:  q   <=  32'b00111110011000000111001101010001 ;
        2690:  q   <=  32'b00111110011000001000010000011000 ;
        2691:  q   <=  32'b00111110011000001001010011011111 ;
        2692:  q   <=  32'b00111110011000001010010110100101 ;
        2693:  q   <=  32'b00111110011000001011011001101010 ;
        2694:  q   <=  32'b00111110011000001100011100101111 ;
        2695:  q   <=  32'b00111110011000001101011111110011 ;
        2696:  q   <=  32'b00111110011000001110100010110110 ;
        2697:  q   <=  32'b00111110011000001111100101111001 ;
        2698:  q   <=  32'b00111110011000010000101000111011 ;
        2699:  q   <=  32'b00111110011000010001101011111100 ;
        2700:  q   <=  32'b00111110011000010010101110111101 ;
        2701:  q   <=  32'b00111110011000010011110001111110 ;
        2702:  q   <=  32'b00111110011000010100110100111101 ;
        2703:  q   <=  32'b00111110011000010101110111111100 ;
        2704:  q   <=  32'b00111110011000010110111010111010 ;
        2705:  q   <=  32'b00111110011000010111111101111000 ;
        2706:  q   <=  32'b00111110011000011001000000110101 ;
        2707:  q   <=  32'b00111110011000011010000011110010 ;
        2708:  q   <=  32'b00111110011000011011000110101110 ;
        2709:  q   <=  32'b00111110011000011100001001101001 ;
        2710:  q   <=  32'b00111110011000011101001100100011 ;
        2711:  q   <=  32'b00111110011000011110001111011101 ;
        2712:  q   <=  32'b00111110011000011111010010010111 ;
        2713:  q   <=  32'b00111110011000100000010101001111 ;
        2714:  q   <=  32'b00111110011000100001011000000111 ;
        2715:  q   <=  32'b00111110011000100010011010111111 ;
        2716:  q   <=  32'b00111110011000100011011101110101 ;
        2717:  q   <=  32'b00111110011000100100100000101100 ;
        2718:  q   <=  32'b00111110011000100101100011100001 ;
        2719:  q   <=  32'b00111110011000100110100110010110 ;
        2720:  q   <=  32'b00111110011000100111101001001010 ;
        2721:  q   <=  32'b00111110011000101000101011111110 ;
        2722:  q   <=  32'b00111110011000101001101110110001 ;
        2723:  q   <=  32'b00111110011000101010110001100011 ;
        2724:  q   <=  32'b00111110011000101011110100010101 ;
        2725:  q   <=  32'b00111110011000101100110111000110 ;
        2726:  q   <=  32'b00111110011000101101111001110111 ;
        2727:  q   <=  32'b00111110011000101110111100100111 ;
        2728:  q   <=  32'b00111110011000101111111111010110 ;
        2729:  q   <=  32'b00111110011000110001000010000101 ;
        2730:  q   <=  32'b00111110011000110010000100110011 ;
        2731:  q   <=  32'b00111110011000110011000111100000 ;
        2732:  q   <=  32'b00111110011000110100001010001101 ;
        2733:  q   <=  32'b00111110011000110101001100111001 ;
        2734:  q   <=  32'b00111110011000110110001111100101 ;
        2735:  q   <=  32'b00111110011000110111010010001111 ;
        2736:  q   <=  32'b00111110011000111000010100111010 ;
        2737:  q   <=  32'b00111110011000111001010111100011 ;
        2738:  q   <=  32'b00111110011000111010011010001100 ;
        2739:  q   <=  32'b00111110011000111011011100110101 ;
        2740:  q   <=  32'b00111110011000111100011111011101 ;
        2741:  q   <=  32'b00111110011000111101100010000100 ;
        2742:  q   <=  32'b00111110011000111110100100101010 ;
        2743:  q   <=  32'b00111110011000111111100111010000 ;
        2744:  q   <=  32'b00111110011001000000101001110101 ;
        2745:  q   <=  32'b00111110011001000001101100011010 ;
        2746:  q   <=  32'b00111110011001000010101110111110 ;
        2747:  q   <=  32'b00111110011001000011110001100001 ;
        2748:  q   <=  32'b00111110011001000100110100000100 ;
        2749:  q   <=  32'b00111110011001000101110110100110 ;
        2750:  q   <=  32'b00111110011001000110111001001000 ;
        2751:  q   <=  32'b00111110011001000111111011101001 ;
        2752:  q   <=  32'b00111110011001001000111110001001 ;
        2753:  q   <=  32'b00111110011001001010000000101001 ;
        2754:  q   <=  32'b00111110011001001011000011001000 ;
        2755:  q   <=  32'b00111110011001001100000101100110 ;
        2756:  q   <=  32'b00111110011001001101001000000100 ;
        2757:  q   <=  32'b00111110011001001110001010100001 ;
        2758:  q   <=  32'b00111110011001001111001100111110 ;
        2759:  q   <=  32'b00111110011001010000001111011010 ;
        2760:  q   <=  32'b00111110011001010001010001110101 ;
        2761:  q   <=  32'b00111110011001010010010100010000 ;
        2762:  q   <=  32'b00111110011001010011010110101010 ;
        2763:  q   <=  32'b00111110011001010100011001000100 ;
        2764:  q   <=  32'b00111110011001010101011011011100 ;
        2765:  q   <=  32'b00111110011001010110011101110101 ;
        2766:  q   <=  32'b00111110011001010111100000001100 ;
        2767:  q   <=  32'b00111110011001011000100010100011 ;
        2768:  q   <=  32'b00111110011001011001100100111010 ;
        2769:  q   <=  32'b00111110011001011010100111001111 ;
        2770:  q   <=  32'b00111110011001011011101001100100 ;
        2771:  q   <=  32'b00111110011001011100101011111001 ;
        2772:  q   <=  32'b00111110011001011101101110001101 ;
        2773:  q   <=  32'b00111110011001011110110000100000 ;
        2774:  q   <=  32'b00111110011001011111110010110011 ;
        2775:  q   <=  32'b00111110011001100000110101000101 ;
        2776:  q   <=  32'b00111110011001100001110111010110 ;
        2777:  q   <=  32'b00111110011001100010111001100111 ;
        2778:  q   <=  32'b00111110011001100011111011110111 ;
        2779:  q   <=  32'b00111110011001100100111110000111 ;
        2780:  q   <=  32'b00111110011001100110000000010110 ;
        2781:  q   <=  32'b00111110011001100111000010100100 ;
        2782:  q   <=  32'b00111110011001101000000100110010 ;
        2783:  q   <=  32'b00111110011001101001000110111111 ;
        2784:  q   <=  32'b00111110011001101010001001001100 ;
        2785:  q   <=  32'b00111110011001101011001011011000 ;
        2786:  q   <=  32'b00111110011001101100001101100011 ;
        2787:  q   <=  32'b00111110011001101101001111101101 ;
        2788:  q   <=  32'b00111110011001101110010001110111 ;
        2789:  q   <=  32'b00111110011001101111010100000001 ;
        2790:  q   <=  32'b00111110011001110000010110001010 ;
        2791:  q   <=  32'b00111110011001110001011000010010 ;
        2792:  q   <=  32'b00111110011001110010011010011001 ;
        2793:  q   <=  32'b00111110011001110011011100100000 ;
        2794:  q   <=  32'b00111110011001110100011110100111 ;
        2795:  q   <=  32'b00111110011001110101100000101101 ;
        2796:  q   <=  32'b00111110011001110110100010110010 ;
        2797:  q   <=  32'b00111110011001110111100100110110 ;
        2798:  q   <=  32'b00111110011001111000100110111010 ;
        2799:  q   <=  32'b00111110011001111001101000111101 ;
        2800:  q   <=  32'b00111110011001111010101011000000 ;
        2801:  q   <=  32'b00111110011001111011101101000010 ;
        2802:  q   <=  32'b00111110011001111100101111000100 ;
        2803:  q   <=  32'b00111110011001111101110001000100 ;
        2804:  q   <=  32'b00111110011001111110110011000101 ;
        2805:  q   <=  32'b00111110011001111111110101000100 ;
        2806:  q   <=  32'b00111110011010000000110111000011 ;
        2807:  q   <=  32'b00111110011010000001111001000010 ;
        2808:  q   <=  32'b00111110011010000010111010111111 ;
        2809:  q   <=  32'b00111110011010000011111100111101 ;
        2810:  q   <=  32'b00111110011010000100111110111001 ;
        2811:  q   <=  32'b00111110011010000110000000110101 ;
        2812:  q   <=  32'b00111110011010000111000010110000 ;
        2813:  q   <=  32'b00111110011010001000000100101011 ;
        2814:  q   <=  32'b00111110011010001001000110100101 ;
        2815:  q   <=  32'b00111110011010001010001000011111 ;
        2816:  q   <=  32'b00111110011010001011001010011000 ;
        2817:  q   <=  32'b00111110011010001100001100010000 ;
        2818:  q   <=  32'b00111110011010001101001110000111 ;
        2819:  q   <=  32'b00111110011010001110001111111111 ;
        2820:  q   <=  32'b00111110011010001111010001110101 ;
        2821:  q   <=  32'b00111110011010010000010011101011 ;
        2822:  q   <=  32'b00111110011010010001010101100000 ;
        2823:  q   <=  32'b00111110011010010010010111010101 ;
        2824:  q   <=  32'b00111110011010010011011001001001 ;
        2825:  q   <=  32'b00111110011010010100011010111100 ;
        2826:  q   <=  32'b00111110011010010101011100101111 ;
        2827:  q   <=  32'b00111110011010010110011110100001 ;
        2828:  q   <=  32'b00111110011010010111100000010011 ;
        2829:  q   <=  32'b00111110011010011000100010000100 ;
        2830:  q   <=  32'b00111110011010011001100011110100 ;
        2831:  q   <=  32'b00111110011010011010100101100100 ;
        2832:  q   <=  32'b00111110011010011011100111010011 ;
        2833:  q   <=  32'b00111110011010011100101001000001 ;
        2834:  q   <=  32'b00111110011010011101101010101111 ;
        2835:  q   <=  32'b00111110011010011110101100011101 ;
        2836:  q   <=  32'b00111110011010011111101110001001 ;
        2837:  q   <=  32'b00111110011010100000101111110101 ;
        2838:  q   <=  32'b00111110011010100001110001100001 ;
        2839:  q   <=  32'b00111110011010100010110011001100 ;
        2840:  q   <=  32'b00111110011010100011110100110110 ;
        2841:  q   <=  32'b00111110011010100100110110100000 ;
        2842:  q   <=  32'b00111110011010100101111000001001 ;
        2843:  q   <=  32'b00111110011010100110111001110001 ;
        2844:  q   <=  32'b00111110011010100111111011011001 ;
        2845:  q   <=  32'b00111110011010101000111101000001 ;
        2846:  q   <=  32'b00111110011010101001111110100111 ;
        2847:  q   <=  32'b00111110011010101011000000001101 ;
        2848:  q   <=  32'b00111110011010101100000001110011 ;
        2849:  q   <=  32'b00111110011010101101000011011000 ;
        2850:  q   <=  32'b00111110011010101110000100111100 ;
        2851:  q   <=  32'b00111110011010101111000110011111 ;
        2852:  q   <=  32'b00111110011010110000001000000011 ;
        2853:  q   <=  32'b00111110011010110001001001100101 ;
        2854:  q   <=  32'b00111110011010110010001011000111 ;
        2855:  q   <=  32'b00111110011010110011001100101000 ;
        2856:  q   <=  32'b00111110011010110100001110001001 ;
        2857:  q   <=  32'b00111110011010110101001111101001 ;
        2858:  q   <=  32'b00111110011010110110010001001000 ;
        2859:  q   <=  32'b00111110011010110111010010100111 ;
        2860:  q   <=  32'b00111110011010111000010100000101 ;
        2861:  q   <=  32'b00111110011010111001010101100011 ;
        2862:  q   <=  32'b00111110011010111010010111000000 ;
        2863:  q   <=  32'b00111110011010111011011000011100 ;
        2864:  q   <=  32'b00111110011010111100011001111000 ;
        2865:  q   <=  32'b00111110011010111101011011010011 ;
        2866:  q   <=  32'b00111110011010111110011100101110 ;
        2867:  q   <=  32'b00111110011010111111011110001000 ;
        2868:  q   <=  32'b00111110011011000000011111100001 ;
        2869:  q   <=  32'b00111110011011000001100000111010 ;
        2870:  q   <=  32'b00111110011011000010100010010010 ;
        2871:  q   <=  32'b00111110011011000011100011101010 ;
        2872:  q   <=  32'b00111110011011000100100101000001 ;
        2873:  q   <=  32'b00111110011011000101100110010111 ;
        2874:  q   <=  32'b00111110011011000110100111101101 ;
        2875:  q   <=  32'b00111110011011000111101001000010 ;
        2876:  q   <=  32'b00111110011011001000101010010111 ;
        2877:  q   <=  32'b00111110011011001001101011101011 ;
        2878:  q   <=  32'b00111110011011001010101100111110 ;
        2879:  q   <=  32'b00111110011011001011101110010001 ;
        2880:  q   <=  32'b00111110011011001100101111100011 ;
        2881:  q   <=  32'b00111110011011001101110000110101 ;
        2882:  q   <=  32'b00111110011011001110110010000110 ;
        2883:  q   <=  32'b00111110011011001111110011010110 ;
        2884:  q   <=  32'b00111110011011010000110100100110 ;
        2885:  q   <=  32'b00111110011011010001110101110101 ;
        2886:  q   <=  32'b00111110011011010010110111000100 ;
        2887:  q   <=  32'b00111110011011010011111000010010 ;
        2888:  q   <=  32'b00111110011011010100111001011111 ;
        2889:  q   <=  32'b00111110011011010101111010101100 ;
        2890:  q   <=  32'b00111110011011010110111011111000 ;
        2891:  q   <=  32'b00111110011011010111111101000100 ;
        2892:  q   <=  32'b00111110011011011000111110001111 ;
        2893:  q   <=  32'b00111110011011011001111111011001 ;
        2894:  q   <=  32'b00111110011011011011000000100011 ;
        2895:  q   <=  32'b00111110011011011100000001101100 ;
        2896:  q   <=  32'b00111110011011011101000010110101 ;
        2897:  q   <=  32'b00111110011011011110000011111101 ;
        2898:  q   <=  32'b00111110011011011111000101000100 ;
        2899:  q   <=  32'b00111110011011100000000110001011 ;
        2900:  q   <=  32'b00111110011011100001000111010001 ;
        2901:  q   <=  32'b00111110011011100010001000010111 ;
        2902:  q   <=  32'b00111110011011100011001001011100 ;
        2903:  q   <=  32'b00111110011011100100001010100001 ;
        2904:  q   <=  32'b00111110011011100101001011100100 ;
        2905:  q   <=  32'b00111110011011100110001100101000 ;
        2906:  q   <=  32'b00111110011011100111001101101010 ;
        2907:  q   <=  32'b00111110011011101000001110101101 ;
        2908:  q   <=  32'b00111110011011101001001111101110 ;
        2909:  q   <=  32'b00111110011011101010010000101111 ;
        2910:  q   <=  32'b00111110011011101011010001101111 ;
        2911:  q   <=  32'b00111110011011101100010010101111 ;
        2912:  q   <=  32'b00111110011011101101010011101110 ;
        2913:  q   <=  32'b00111110011011101110010100101101 ;
        2914:  q   <=  32'b00111110011011101111010101101010 ;
        2915:  q   <=  32'b00111110011011110000010110101000 ;
        2916:  q   <=  32'b00111110011011110001010111100101 ;
        2917:  q   <=  32'b00111110011011110010011000100001 ;
        2918:  q   <=  32'b00111110011011110011011001011100 ;
        2919:  q   <=  32'b00111110011011110100011010010111 ;
        2920:  q   <=  32'b00111110011011110101011011010010 ;
        2921:  q   <=  32'b00111110011011110110011100001011 ;
        2922:  q   <=  32'b00111110011011110111011101000101 ;
        2923:  q   <=  32'b00111110011011111000011101111101 ;
        2924:  q   <=  32'b00111110011011111001011110110101 ;
        2925:  q   <=  32'b00111110011011111010011111101101 ;
        2926:  q   <=  32'b00111110011011111011100000100011 ;
        2927:  q   <=  32'b00111110011011111100100001011010 ;
        2928:  q   <=  32'b00111110011011111101100010001111 ;
        2929:  q   <=  32'b00111110011011111110100011000100 ;
        2930:  q   <=  32'b00111110011011111111100011111001 ;
        2931:  q   <=  32'b00111110011100000000100100101101 ;
        2932:  q   <=  32'b00111110011100000001100101100000 ;
        2933:  q   <=  32'b00111110011100000010100110010011 ;
        2934:  q   <=  32'b00111110011100000011100111000101 ;
        2935:  q   <=  32'b00111110011100000100100111110110 ;
        2936:  q   <=  32'b00111110011100000101101000100111 ;
        2937:  q   <=  32'b00111110011100000110101001011000 ;
        2938:  q   <=  32'b00111110011100000111101010000111 ;
        2939:  q   <=  32'b00111110011100001000101010110110 ;
        2940:  q   <=  32'b00111110011100001001101011100101 ;
        2941:  q   <=  32'b00111110011100001010101100010011 ;
        2942:  q   <=  32'b00111110011100001011101101000000 ;
        2943:  q   <=  32'b00111110011100001100101101101101 ;
        2944:  q   <=  32'b00111110011100001101101110011001 ;
        2945:  q   <=  32'b00111110011100001110101111000101 ;
        2946:  q   <=  32'b00111110011100001111101111110000 ;
        2947:  q   <=  32'b00111110011100010000110000011010 ;
        2948:  q   <=  32'b00111110011100010001110001000100 ;
        2949:  q   <=  32'b00111110011100010010110001101110 ;
        2950:  q   <=  32'b00111110011100010011110010010110 ;
        2951:  q   <=  32'b00111110011100010100110010111110 ;
        2952:  q   <=  32'b00111110011100010101110011100110 ;
        2953:  q   <=  32'b00111110011100010110110100001101 ;
        2954:  q   <=  32'b00111110011100010111110100110011 ;
        2955:  q   <=  32'b00111110011100011000110101011001 ;
        2956:  q   <=  32'b00111110011100011001110101111110 ;
        2957:  q   <=  32'b00111110011100011010110110100011 ;
        2958:  q   <=  32'b00111110011100011011110111000111 ;
        2959:  q   <=  32'b00111110011100011100110111101010 ;
        2960:  q   <=  32'b00111110011100011101111000001101 ;
        2961:  q   <=  32'b00111110011100011110111000101111 ;
        2962:  q   <=  32'b00111110011100011111111001010001 ;
        2963:  q   <=  32'b00111110011100100000111001110010 ;
        2964:  q   <=  32'b00111110011100100001111010010010 ;
        2965:  q   <=  32'b00111110011100100010111010110010 ;
        2966:  q   <=  32'b00111110011100100011111011010001 ;
        2967:  q   <=  32'b00111110011100100100111011110000 ;
        2968:  q   <=  32'b00111110011100100101111100001110 ;
        2969:  q   <=  32'b00111110011100100110111100101100 ;
        2970:  q   <=  32'b00111110011100100111111101001001 ;
        2971:  q   <=  32'b00111110011100101000111101100101 ;
        2972:  q   <=  32'b00111110011100101001111110000001 ;
        2973:  q   <=  32'b00111110011100101010111110011100 ;
        2974:  q   <=  32'b00111110011100101011111110110111 ;
        2975:  q   <=  32'b00111110011100101100111111010001 ;
        2976:  q   <=  32'b00111110011100101101111111101010 ;
        2977:  q   <=  32'b00111110011100101111000000000011 ;
        2978:  q   <=  32'b00111110011100110000000000011100 ;
        2979:  q   <=  32'b00111110011100110001000000110011 ;
        2980:  q   <=  32'b00111110011100110010000001001011 ;
        2981:  q   <=  32'b00111110011100110011000001100001 ;
        2982:  q   <=  32'b00111110011100110100000001110111 ;
        2983:  q   <=  32'b00111110011100110101000010001101 ;
        2984:  q   <=  32'b00111110011100110110000010100001 ;
        2985:  q   <=  32'b00111110011100110111000010110110 ;
        2986:  q   <=  32'b00111110011100111000000011001001 ;
        2987:  q   <=  32'b00111110011100111001000011011100 ;
        2988:  q   <=  32'b00111110011100111010000011101111 ;
        2989:  q   <=  32'b00111110011100111011000100000001 ;
        2990:  q   <=  32'b00111110011100111100000100010010 ;
        2991:  q   <=  32'b00111110011100111101000100100011 ;
        2992:  q   <=  32'b00111110011100111110000100110011 ;
        2993:  q   <=  32'b00111110011100111111000101000011 ;
        2994:  q   <=  32'b00111110011101000000000101010010 ;
        2995:  q   <=  32'b00111110011101000001000101100000 ;
        2996:  q   <=  32'b00111110011101000010000101101110 ;
        2997:  q   <=  32'b00111110011101000011000101111011 ;
        2998:  q   <=  32'b00111110011101000100000110001000 ;
        2999:  q   <=  32'b00111110011101000101000110010100 ;
        3000:  q   <=  32'b00111110011101000110000110011111 ;
        3001:  q   <=  32'b00111110011101000111000110101010 ;
        3002:  q   <=  32'b00111110011101001000000110110101 ;
        3003:  q   <=  32'b00111110011101001001000110111111 ;
        3004:  q   <=  32'b00111110011101001010000111001000 ;
        3005:  q   <=  32'b00111110011101001011000111010000 ;
        3006:  q   <=  32'b00111110011101001100000111011000 ;
        3007:  q   <=  32'b00111110011101001101000111100000 ;
        3008:  q   <=  32'b00111110011101001110000111100111 ;
        3009:  q   <=  32'b00111110011101001111000111101101 ;
        3010:  q   <=  32'b00111110011101010000000111110011 ;
        3011:  q   <=  32'b00111110011101010001000111111000 ;
        3012:  q   <=  32'b00111110011101010010000111111101 ;
        3013:  q   <=  32'b00111110011101010011001000000001 ;
        3014:  q   <=  32'b00111110011101010100001000000100 ;
        3015:  q   <=  32'b00111110011101010101001000000111 ;
        3016:  q   <=  32'b00111110011101010110001000001001 ;
        3017:  q   <=  32'b00111110011101010111001000001011 ;
        3018:  q   <=  32'b00111110011101011000001000001100 ;
        3019:  q   <=  32'b00111110011101011001001000001101 ;
        3020:  q   <=  32'b00111110011101011010001000001101 ;
        3021:  q   <=  32'b00111110011101011011001000001100 ;
        3022:  q   <=  32'b00111110011101011100001000001011 ;
        3023:  q   <=  32'b00111110011101011101001000001001 ;
        3024:  q   <=  32'b00111110011101011110001000000111 ;
        3025:  q   <=  32'b00111110011101011111001000000100 ;
        3026:  q   <=  32'b00111110011101100000001000000001 ;
        3027:  q   <=  32'b00111110011101100001000111111101 ;
        3028:  q   <=  32'b00111110011101100010000111111000 ;
        3029:  q   <=  32'b00111110011101100011000111110011 ;
        3030:  q   <=  32'b00111110011101100100000111101101 ;
        3031:  q   <=  32'b00111110011101100101000111100111 ;
        3032:  q   <=  32'b00111110011101100110000111100000 ;
        3033:  q   <=  32'b00111110011101100111000111011000 ;
        3034:  q   <=  32'b00111110011101101000000111010000 ;
        3035:  q   <=  32'b00111110011101101001000111001000 ;
        3036:  q   <=  32'b00111110011101101010000110111110 ;
        3037:  q   <=  32'b00111110011101101011000110110101 ;
        3038:  q   <=  32'b00111110011101101100000110101010 ;
        3039:  q   <=  32'b00111110011101101101000110011111 ;
        3040:  q   <=  32'b00111110011101101110000110010100 ;
        3041:  q   <=  32'b00111110011101101111000110001000 ;
        3042:  q   <=  32'b00111110011101110000000101111011 ;
        3043:  q   <=  32'b00111110011101110001000101101110 ;
        3044:  q   <=  32'b00111110011101110010000101100000 ;
        3045:  q   <=  32'b00111110011101110011000101010010 ;
        3046:  q   <=  32'b00111110011101110100000101000011 ;
        3047:  q   <=  32'b00111110011101110101000100110011 ;
        3048:  q   <=  32'b00111110011101110110000100100011 ;
        3049:  q   <=  32'b00111110011101110111000100010011 ;
        3050:  q   <=  32'b00111110011101111000000100000010 ;
        3051:  q   <=  32'b00111110011101111001000011110000 ;
        3052:  q   <=  32'b00111110011101111010000011011101 ;
        3053:  q   <=  32'b00111110011101111011000011001010 ;
        3054:  q   <=  32'b00111110011101111100000010110111 ;
        3055:  q   <=  32'b00111110011101111101000010100011 ;
        3056:  q   <=  32'b00111110011101111110000010001110 ;
        3057:  q   <=  32'b00111110011101111111000001111001 ;
        3058:  q   <=  32'b00111110011110000000000001100011 ;
        3059:  q   <=  32'b00111110011110000001000001001101 ;
        3060:  q   <=  32'b00111110011110000010000000110110 ;
        3061:  q   <=  32'b00111110011110000011000000011111 ;
        3062:  q   <=  32'b00111110011110000100000000000111 ;
        3063:  q   <=  32'b00111110011110000100111111101110 ;
        3064:  q   <=  32'b00111110011110000101111111010101 ;
        3065:  q   <=  32'b00111110011110000110111110111011 ;
        3066:  q   <=  32'b00111110011110000111111110100001 ;
        3067:  q   <=  32'b00111110011110001000111110000110 ;
        3068:  q   <=  32'b00111110011110001001111101101010 ;
        3069:  q   <=  32'b00111110011110001010111101001110 ;
        3070:  q   <=  32'b00111110011110001011111100110010 ;
        3071:  q   <=  32'b00111110011110001100111100010101 ;
        3072:  q   <=  32'b00111110011110001101111011110111 ;
        3073:  q   <=  32'b00111110011110001110111011011001 ;
        3074:  q   <=  32'b00111110011110001111111010111010 ;
        3075:  q   <=  32'b00111110011110010000111010011010 ;
        3076:  q   <=  32'b00111110011110010001111001111010 ;
        3077:  q   <=  32'b00111110011110010010111001011010 ;
        3078:  q   <=  32'b00111110011110010011111000111001 ;
        3079:  q   <=  32'b00111110011110010100111000010111 ;
        3080:  q   <=  32'b00111110011110010101110111110101 ;
        3081:  q   <=  32'b00111110011110010110110111010010 ;
        3082:  q   <=  32'b00111110011110010111110110101110 ;
        3083:  q   <=  32'b00111110011110011000110110001010 ;
        3084:  q   <=  32'b00111110011110011001110101100110 ;
        3085:  q   <=  32'b00111110011110011010110101000001 ;
        3086:  q   <=  32'b00111110011110011011110100011011 ;
        3087:  q   <=  32'b00111110011110011100110011110101 ;
        3088:  q   <=  32'b00111110011110011101110011001110 ;
        3089:  q   <=  32'b00111110011110011110110010100111 ;
        3090:  q   <=  32'b00111110011110011111110001111111 ;
        3091:  q   <=  32'b00111110011110100000110001010110 ;
        3092:  q   <=  32'b00111110011110100001110000101101 ;
        3093:  q   <=  32'b00111110011110100010110000000100 ;
        3094:  q   <=  32'b00111110011110100011101111011010 ;
        3095:  q   <=  32'b00111110011110100100101110101111 ;
        3096:  q   <=  32'b00111110011110100101101110000100 ;
        3097:  q   <=  32'b00111110011110100110101101011000 ;
        3098:  q   <=  32'b00111110011110100111101100101011 ;
        3099:  q   <=  32'b00111110011110101000101011111110 ;
        3100:  q   <=  32'b00111110011110101001101011010001 ;
        3101:  q   <=  32'b00111110011110101010101010100011 ;
        3102:  q   <=  32'b00111110011110101011101001110100 ;
        3103:  q   <=  32'b00111110011110101100101001000101 ;
        3104:  q   <=  32'b00111110011110101101101000010101 ;
        3105:  q   <=  32'b00111110011110101110100111100101 ;
        3106:  q   <=  32'b00111110011110101111100110110100 ;
        3107:  q   <=  32'b00111110011110110000100110000010 ;
        3108:  q   <=  32'b00111110011110110001100101010000 ;
        3109:  q   <=  32'b00111110011110110010100100011110 ;
        3110:  q   <=  32'b00111110011110110011100011101010 ;
        3111:  q   <=  32'b00111110011110110100100010110111 ;
        3112:  q   <=  32'b00111110011110110101100010000010 ;
        3113:  q   <=  32'b00111110011110110110100001001101 ;
        3114:  q   <=  32'b00111110011110110111100000011000 ;
        3115:  q   <=  32'b00111110011110111000011111100010 ;
        3116:  q   <=  32'b00111110011110111001011110101100 ;
        3117:  q   <=  32'b00111110011110111010011101110100 ;
        3118:  q   <=  32'b00111110011110111011011100111101 ;
        3119:  q   <=  32'b00111110011110111100011100000101 ;
        3120:  q   <=  32'b00111110011110111101011011001100 ;
        3121:  q   <=  32'b00111110011110111110011010010010 ;
        3122:  q   <=  32'b00111110011110111111011001011001 ;
        3123:  q   <=  32'b00111110011111000000011000011110 ;
        3124:  q   <=  32'b00111110011111000001010111100011 ;
        3125:  q   <=  32'b00111110011111000010010110100111 ;
        3126:  q   <=  32'b00111110011111000011010101101011 ;
        3127:  q   <=  32'b00111110011111000100010100101111 ;
        3128:  q   <=  32'b00111110011111000101010011110001 ;
        3129:  q   <=  32'b00111110011111000110010010110100 ;
        3130:  q   <=  32'b00111110011111000111010001110101 ;
        3131:  q   <=  32'b00111110011111001000010000110110 ;
        3132:  q   <=  32'b00111110011111001001001111110111 ;
        3133:  q   <=  32'b00111110011111001010001110110111 ;
        3134:  q   <=  32'b00111110011111001011001101110110 ;
        3135:  q   <=  32'b00111110011111001100001100110101 ;
        3136:  q   <=  32'b00111110011111001101001011110011 ;
        3137:  q   <=  32'b00111110011111001110001010110001 ;
        3138:  q   <=  32'b00111110011111001111001001101110 ;
        3139:  q   <=  32'b00111110011111010000001000101011 ;
        3140:  q   <=  32'b00111110011111010001000111100111 ;
        3141:  q   <=  32'b00111110011111010010000110100010 ;
        3142:  q   <=  32'b00111110011111010011000101011101 ;
        3143:  q   <=  32'b00111110011111010100000100011000 ;
        3144:  q   <=  32'b00111110011111010101000011010010 ;
        3145:  q   <=  32'b00111110011111010110000010001011 ;
        3146:  q   <=  32'b00111110011111010111000001000100 ;
        3147:  q   <=  32'b00111110011111010111111111111100 ;
        3148:  q   <=  32'b00111110011111011000111110110011 ;
        3149:  q   <=  32'b00111110011111011001111101101010 ;
        3150:  q   <=  32'b00111110011111011010111100100001 ;
        3151:  q   <=  32'b00111110011111011011111011010111 ;
        3152:  q   <=  32'b00111110011111011100111010001100 ;
        3153:  q   <=  32'b00111110011111011101111001000001 ;
        3154:  q   <=  32'b00111110011111011110110111110101 ;
        3155:  q   <=  32'b00111110011111011111110110101001 ;
        3156:  q   <=  32'b00111110011111100000110101011100 ;
        3157:  q   <=  32'b00111110011111100001110100001111 ;
        3158:  q   <=  32'b00111110011111100010110011000001 ;
        3159:  q   <=  32'b00111110011111100011110001110010 ;
        3160:  q   <=  32'b00111110011111100100110000100011 ;
        3161:  q   <=  32'b00111110011111100101101111010100 ;
        3162:  q   <=  32'b00111110011111100110101110000100 ;
        3163:  q   <=  32'b00111110011111100111101100110011 ;
        3164:  q   <=  32'b00111110011111101000101011100010 ;
        3165:  q   <=  32'b00111110011111101001101010010000 ;
        3166:  q   <=  32'b00111110011111101010101000111101 ;
        3167:  q   <=  32'b00111110011111101011100111101011 ;
        3168:  q   <=  32'b00111110011111101100100110010111 ;
        3169:  q   <=  32'b00111110011111101101100101000011 ;
        3170:  q   <=  32'b00111110011111101110100011101110 ;
        3171:  q   <=  32'b00111110011111101111100010011001 ;
        3172:  q   <=  32'b00111110011111110000100001000100 ;
        3173:  q   <=  32'b00111110011111110001011111101101 ;
        3174:  q   <=  32'b00111110011111110010011110010111 ;
        3175:  q   <=  32'b00111110011111110011011100111111 ;
        3176:  q   <=  32'b00111110011111110100011011100111 ;
        3177:  q   <=  32'b00111110011111110101011010001111 ;
        3178:  q   <=  32'b00111110011111110110011000110110 ;
        3179:  q   <=  32'b00111110011111110111010111011100 ;
        3180:  q   <=  32'b00111110011111111000010110000010 ;
        3181:  q   <=  32'b00111110011111111001010100101000 ;
        3182:  q   <=  32'b00111110011111111010010011001101 ;
        3183:  q   <=  32'b00111110011111111011010001110001 ;
        3184:  q   <=  32'b00111110011111111100010000010101 ;
        3185:  q   <=  32'b00111110011111111101001110111000 ;
        3186:  q   <=  32'b00111110011111111110001101011010 ;
        3187:  q   <=  32'b00111110011111111111001011111100 ;
        3188:  q   <=  32'b00111110100000000000000101001111 ;
        3189:  q   <=  32'b00111110100000000000100100011111 ;
        3190:  q   <=  32'b00111110100000000001000011101111 ;
        3191:  q   <=  32'b00111110100000000001100010111111 ;
        3192:  q   <=  32'b00111110100000000010000010001111 ;
        3193:  q   <=  32'b00111110100000000010100001011110 ;
        3194:  q   <=  32'b00111110100000000011000000101101 ;
        3195:  q   <=  32'b00111110100000000011011111111100 ;
        3196:  q   <=  32'b00111110100000000011111111001011 ;
        3197:  q   <=  32'b00111110100000000100011110011001 ;
        3198:  q   <=  32'b00111110100000000100111101100111 ;
        3199:  q   <=  32'b00111110100000000101011100110101 ;
        3200:  q   <=  32'b00111110100000000101111100000010 ;
        3201:  q   <=  32'b00111110100000000110011011010000 ;
        3202:  q   <=  32'b00111110100000000110111010011100 ;
        3203:  q   <=  32'b00111110100000000111011001101001 ;
        3204:  q   <=  32'b00111110100000000111111000110101 ;
        3205:  q   <=  32'b00111110100000001000011000000010 ;
        3206:  q   <=  32'b00111110100000001000110111001101 ;
        3207:  q   <=  32'b00111110100000001001010110011001 ;
        3208:  q   <=  32'b00111110100000001001110101100100 ;
        3209:  q   <=  32'b00111110100000001010010100101111 ;
        3210:  q   <=  32'b00111110100000001010110011111010 ;
        3211:  q   <=  32'b00111110100000001011010011000100 ;
        3212:  q   <=  32'b00111110100000001011110010001111 ;
        3213:  q   <=  32'b00111110100000001100010001011001 ;
        3214:  q   <=  32'b00111110100000001100110000100010 ;
        3215:  q   <=  32'b00111110100000001101001111101100 ;
        3216:  q   <=  32'b00111110100000001101101110110101 ;
        3217:  q   <=  32'b00111110100000001110001101111101 ;
        3218:  q   <=  32'b00111110100000001110101101000110 ;
        3219:  q   <=  32'b00111110100000001111001100001110 ;
        3220:  q   <=  32'b00111110100000001111101011010110 ;
        3221:  q   <=  32'b00111110100000010000001010011110 ;
        3222:  q   <=  32'b00111110100000010000101001100101 ;
        3223:  q   <=  32'b00111110100000010001001000101101 ;
        3224:  q   <=  32'b00111110100000010001100111110100 ;
        3225:  q   <=  32'b00111110100000010010000110111010 ;
        3226:  q   <=  32'b00111110100000010010100110000001 ;
        3227:  q   <=  32'b00111110100000010011000101000111 ;
        3228:  q   <=  32'b00111110100000010011100100001100 ;
        3229:  q   <=  32'b00111110100000010100000011010010 ;
        3230:  q   <=  32'b00111110100000010100100010010111 ;
        3231:  q   <=  32'b00111110100000010101000001011100 ;
        3232:  q   <=  32'b00111110100000010101100000100001 ;
        3233:  q   <=  32'b00111110100000010101111111100110 ;
        3234:  q   <=  32'b00111110100000010110011110101010 ;
        3235:  q   <=  32'b00111110100000010110111101101110 ;
        3236:  q   <=  32'b00111110100000010111011100110001 ;
        3237:  q   <=  32'b00111110100000010111111011110101 ;
        3238:  q   <=  32'b00111110100000011000011010111000 ;
        3239:  q   <=  32'b00111110100000011000111001111011 ;
        3240:  q   <=  32'b00111110100000011001011000111101 ;
        3241:  q   <=  32'b00111110100000011001111000000000 ;
        3242:  q   <=  32'b00111110100000011010010111000010 ;
        3243:  q   <=  32'b00111110100000011010110110000011 ;
        3244:  q   <=  32'b00111110100000011011010101000101 ;
        3245:  q   <=  32'b00111110100000011011110100000110 ;
        3246:  q   <=  32'b00111110100000011100010011000111 ;
        3247:  q   <=  32'b00111110100000011100110010001000 ;
        3248:  q   <=  32'b00111110100000011101010001001000 ;
        3249:  q   <=  32'b00111110100000011101110000001000 ;
        3250:  q   <=  32'b00111110100000011110001111001000 ;
        3251:  q   <=  32'b00111110100000011110101110001000 ;
        3252:  q   <=  32'b00111110100000011111001101000111 ;
        3253:  q   <=  32'b00111110100000011111101100000110 ;
        3254:  q   <=  32'b00111110100000100000001011000101 ;
        3255:  q   <=  32'b00111110100000100000101010000011 ;
        3256:  q   <=  32'b00111110100000100001001001000010 ;
        3257:  q   <=  32'b00111110100000100001101000000000 ;
        3258:  q   <=  32'b00111110100000100010000110111101 ;
        3259:  q   <=  32'b00111110100000100010100101111011 ;
        3260:  q   <=  32'b00111110100000100011000100111000 ;
        3261:  q   <=  32'b00111110100000100011100011110101 ;
        3262:  q   <=  32'b00111110100000100100000010110001 ;
        3263:  q   <=  32'b00111110100000100100100001101110 ;
        3264:  q   <=  32'b00111110100000100101000000101010 ;
        3265:  q   <=  32'b00111110100000100101011111100110 ;
        3266:  q   <=  32'b00111110100000100101111110100001 ;
        3267:  q   <=  32'b00111110100000100110011101011101 ;
        3268:  q   <=  32'b00111110100000100110111100011000 ;
        3269:  q   <=  32'b00111110100000100111011011010010 ;
        3270:  q   <=  32'b00111110100000100111111010001101 ;
        3271:  q   <=  32'b00111110100000101000011001000111 ;
        3272:  q   <=  32'b00111110100000101000111000000001 ;
        3273:  q   <=  32'b00111110100000101001010110111011 ;
        3274:  q   <=  32'b00111110100000101001110101110100 ;
        3275:  q   <=  32'b00111110100000101010010100101101 ;
        3276:  q   <=  32'b00111110100000101010110011100110 ;
        3277:  q   <=  32'b00111110100000101011010010011111 ;
        3278:  q   <=  32'b00111110100000101011110001010111 ;
        3279:  q   <=  32'b00111110100000101100010000001111 ;
        3280:  q   <=  32'b00111110100000101100101111000111 ;
        3281:  q   <=  32'b00111110100000101101001101111110 ;
        3282:  q   <=  32'b00111110100000101101101100110110 ;
        3283:  q   <=  32'b00111110100000101110001011101101 ;
        3284:  q   <=  32'b00111110100000101110101010100011 ;
        3285:  q   <=  32'b00111110100000101111001001011010 ;
        3286:  q   <=  32'b00111110100000101111101000010000 ;
        3287:  q   <=  32'b00111110100000110000000111000110 ;
        3288:  q   <=  32'b00111110100000110000100101111100 ;
        3289:  q   <=  32'b00111110100000110001000100110001 ;
        3290:  q   <=  32'b00111110100000110001100011100110 ;
        3291:  q   <=  32'b00111110100000110010000010011011 ;
        3292:  q   <=  32'b00111110100000110010100001010000 ;
        3293:  q   <=  32'b00111110100000110011000000000100 ;
        3294:  q   <=  32'b00111110100000110011011110111000 ;
        3295:  q   <=  32'b00111110100000110011111101101100 ;
        3296:  q   <=  32'b00111110100000110100011100011111 ;
        3297:  q   <=  32'b00111110100000110100111011010011 ;
        3298:  q   <=  32'b00111110100000110101011010000110 ;
        3299:  q   <=  32'b00111110100000110101111000111000 ;
        3300:  q   <=  32'b00111110100000110110010111101011 ;
        3301:  q   <=  32'b00111110100000110110110110011101 ;
        3302:  q   <=  32'b00111110100000110111010101001111 ;
        3303:  q   <=  32'b00111110100000110111110100000001 ;
        3304:  q   <=  32'b00111110100000111000010010110010 ;
        3305:  q   <=  32'b00111110100000111000110001100011 ;
        3306:  q   <=  32'b00111110100000111001010000010100 ;
        3307:  q   <=  32'b00111110100000111001101111000100 ;
        3308:  q   <=  32'b00111110100000111010001101110101 ;
        3309:  q   <=  32'b00111110100000111010101100100101 ;
        3310:  q   <=  32'b00111110100000111011001011010101 ;
        3311:  q   <=  32'b00111110100000111011101010000100 ;
        3312:  q   <=  32'b00111110100000111100001000110011 ;
        3313:  q   <=  32'b00111110100000111100100111100010 ;
        3314:  q   <=  32'b00111110100000111101000110010001 ;
        3315:  q   <=  32'b00111110100000111101100101000000 ;
        3316:  q   <=  32'b00111110100000111110000011101110 ;
        3317:  q   <=  32'b00111110100000111110100010011100 ;
        3318:  q   <=  32'b00111110100000111111000001001001 ;
        3319:  q   <=  32'b00111110100000111111011111110111 ;
        3320:  q   <=  32'b00111110100000111111111110100100 ;
        3321:  q   <=  32'b00111110100001000000011101010001 ;
        3322:  q   <=  32'b00111110100001000000111011111101 ;
        3323:  q   <=  32'b00111110100001000001011010101010 ;
        3324:  q   <=  32'b00111110100001000001111001010110 ;
        3325:  q   <=  32'b00111110100001000010011000000010 ;
        3326:  q   <=  32'b00111110100001000010110110101101 ;
        3327:  q   <=  32'b00111110100001000011010101011001 ;
        3328:  q   <=  32'b00111110100001000011110100000100 ;
        3329:  q   <=  32'b00111110100001000100010010101110 ;
        3330:  q   <=  32'b00111110100001000100110001011001 ;
        3331:  q   <=  32'b00111110100001000101010000000011 ;
        3332:  q   <=  32'b00111110100001000101101110101101 ;
        3333:  q   <=  32'b00111110100001000110001101010111 ;
        3334:  q   <=  32'b00111110100001000110101100000000 ;
        3335:  q   <=  32'b00111110100001000111001010101001 ;
        3336:  q   <=  32'b00111110100001000111101001010010 ;
        3337:  q   <=  32'b00111110100001001000000111111011 ;
        3338:  q   <=  32'b00111110100001001000100110100011 ;
        3339:  q   <=  32'b00111110100001001001000101001011 ;
        3340:  q   <=  32'b00111110100001001001100011110011 ;
        3341:  q   <=  32'b00111110100001001010000010011011 ;
        3342:  q   <=  32'b00111110100001001010100001000010 ;
        3343:  q   <=  32'b00111110100001001010111111101001 ;
        3344:  q   <=  32'b00111110100001001011011110010000 ;
        3345:  q   <=  32'b00111110100001001011111100110111 ;
        3346:  q   <=  32'b00111110100001001100011011011101 ;
        3347:  q   <=  32'b00111110100001001100111010000011 ;
        3348:  q   <=  32'b00111110100001001101011000101001 ;
        3349:  q   <=  32'b00111110100001001101110111001110 ;
        3350:  q   <=  32'b00111110100001001110010101110011 ;
        3351:  q   <=  32'b00111110100001001110110100011000 ;
        3352:  q   <=  32'b00111110100001001111010010111101 ;
        3353:  q   <=  32'b00111110100001001111110001100001 ;
        3354:  q   <=  32'b00111110100001010000010000000110 ;
        3355:  q   <=  32'b00111110100001010000101110101010 ;
        3356:  q   <=  32'b00111110100001010001001101001101 ;
        3357:  q   <=  32'b00111110100001010001101011110001 ;
        3358:  q   <=  32'b00111110100001010010001010010100 ;
        3359:  q   <=  32'b00111110100001010010101000110111 ;
        3360:  q   <=  32'b00111110100001010011000111011001 ;
        3361:  q   <=  32'b00111110100001010011100101111011 ;
        3362:  q   <=  32'b00111110100001010100000100011110 ;
        3363:  q   <=  32'b00111110100001010100100010111111 ;
        3364:  q   <=  32'b00111110100001010101000001100001 ;
        3365:  q   <=  32'b00111110100001010101100000000010 ;
        3366:  q   <=  32'b00111110100001010101111110100011 ;
        3367:  q   <=  32'b00111110100001010110011101000100 ;
        3368:  q   <=  32'b00111110100001010110111011100100 ;
        3369:  q   <=  32'b00111110100001010111011010000101 ;
        3370:  q   <=  32'b00111110100001010111111000100101 ;
        3371:  q   <=  32'b00111110100001011000010111000100 ;
        3372:  q   <=  32'b00111110100001011000110101100100 ;
        3373:  q   <=  32'b00111110100001011001010100000011 ;
        3374:  q   <=  32'b00111110100001011001110010100010 ;
        3375:  q   <=  32'b00111110100001011010010001000001 ;
        3376:  q   <=  32'b00111110100001011010101111011111 ;
        3377:  q   <=  32'b00111110100001011011001101111101 ;
        3378:  q   <=  32'b00111110100001011011101100011011 ;
        3379:  q   <=  32'b00111110100001011100001010111001 ;
        3380:  q   <=  32'b00111110100001011100101001010110 ;
        3381:  q   <=  32'b00111110100001011101000111110011 ;
        3382:  q   <=  32'b00111110100001011101100110010000 ;
        3383:  q   <=  32'b00111110100001011110000100101101 ;
        3384:  q   <=  32'b00111110100001011110100011001001 ;
        3385:  q   <=  32'b00111110100001011111000001100101 ;
        3386:  q   <=  32'b00111110100001011111100000000001 ;
        3387:  q   <=  32'b00111110100001011111111110011100 ;
        3388:  q   <=  32'b00111110100001100000011100111000 ;
        3389:  q   <=  32'b00111110100001100000111011010011 ;
        3390:  q   <=  32'b00111110100001100001011001101101 ;
        3391:  q   <=  32'b00111110100001100001111000001000 ;
        3392:  q   <=  32'b00111110100001100010010110100010 ;
        3393:  q   <=  32'b00111110100001100010110100111100 ;
        3394:  q   <=  32'b00111110100001100011010011010110 ;
        3395:  q   <=  32'b00111110100001100011110001101111 ;
        3396:  q   <=  32'b00111110100001100100010000001001 ;
        3397:  q   <=  32'b00111110100001100100101110100010 ;
        3398:  q   <=  32'b00111110100001100101001100111010 ;
        3399:  q   <=  32'b00111110100001100101101011010011 ;
        3400:  q   <=  32'b00111110100001100110001001101011 ;
        3401:  q   <=  32'b00111110100001100110101000000011 ;
        3402:  q   <=  32'b00111110100001100111000110011010 ;
        3403:  q   <=  32'b00111110100001100111100100110010 ;
        3404:  q   <=  32'b00111110100001101000000011001001 ;
        3405:  q   <=  32'b00111110100001101000100001100000 ;
        3406:  q   <=  32'b00111110100001101000111111110110 ;
        3407:  q   <=  32'b00111110100001101001011110001101 ;
        3408:  q   <=  32'b00111110100001101001111100100011 ;
        3409:  q   <=  32'b00111110100001101010011010111001 ;
        3410:  q   <=  32'b00111110100001101010111001001110 ;
        3411:  q   <=  32'b00111110100001101011010111100100 ;
        3412:  q   <=  32'b00111110100001101011110101111001 ;
        3413:  q   <=  32'b00111110100001101100010100001101 ;
        3414:  q   <=  32'b00111110100001101100110010100010 ;
        3415:  q   <=  32'b00111110100001101101010000110110 ;
        3416:  q   <=  32'b00111110100001101101101111001010 ;
        3417:  q   <=  32'b00111110100001101110001101011110 ;
        3418:  q   <=  32'b00111110100001101110101011110010 ;
        3419:  q   <=  32'b00111110100001101111001010000101 ;
        3420:  q   <=  32'b00111110100001101111101000011000 ;
        3421:  q   <=  32'b00111110100001110000000110101011 ;
        3422:  q   <=  32'b00111110100001110000100100111101 ;
        3423:  q   <=  32'b00111110100001110001000011001111 ;
        3424:  q   <=  32'b00111110100001110001100001100001 ;
        3425:  q   <=  32'b00111110100001110001111111110011 ;
        3426:  q   <=  32'b00111110100001110010011110000100 ;
        3427:  q   <=  32'b00111110100001110010111100010110 ;
        3428:  q   <=  32'b00111110100001110011011010100110 ;
        3429:  q   <=  32'b00111110100001110011111000110111 ;
        3430:  q   <=  32'b00111110100001110100010111001000 ;
        3431:  q   <=  32'b00111110100001110100110101011000 ;
        3432:  q   <=  32'b00111110100001110101010011101000 ;
        3433:  q   <=  32'b00111110100001110101110001110111 ;
        3434:  q   <=  32'b00111110100001110110010000000111 ;
        3435:  q   <=  32'b00111110100001110110101110010110 ;
        3436:  q   <=  32'b00111110100001110111001100100101 ;
        3437:  q   <=  32'b00111110100001110111101010110011 ;
        3438:  q   <=  32'b00111110100001111000001001000010 ;
        3439:  q   <=  32'b00111110100001111000100111010000 ;
        3440:  q   <=  32'b00111110100001111001000101011110 ;
        3441:  q   <=  32'b00111110100001111001100011101011 ;
        3442:  q   <=  32'b00111110100001111010000001111001 ;
        3443:  q   <=  32'b00111110100001111010100000000110 ;
        3444:  q   <=  32'b00111110100001111010111110010010 ;
        3445:  q   <=  32'b00111110100001111011011100011111 ;
        3446:  q   <=  32'b00111110100001111011111010101011 ;
        3447:  q   <=  32'b00111110100001111100011000110111 ;
        3448:  q   <=  32'b00111110100001111100110111000011 ;
        3449:  q   <=  32'b00111110100001111101010101001111 ;
        3450:  q   <=  32'b00111110100001111101110011011010 ;
        3451:  q   <=  32'b00111110100001111110010001100101 ;
        3452:  q   <=  32'b00111110100001111110101111110000 ;
        3453:  q   <=  32'b00111110100001111111001101111010 ;
        3454:  q   <=  32'b00111110100001111111101100000101 ;
        3455:  q   <=  32'b00111110100010000000001010001111 ;
        3456:  q   <=  32'b00111110100010000000101000011000 ;
        3457:  q   <=  32'b00111110100010000001000110100010 ;
        3458:  q   <=  32'b00111110100010000001100100101011 ;
        3459:  q   <=  32'b00111110100010000010000010110100 ;
        3460:  q   <=  32'b00111110100010000010100000111101 ;
        3461:  q   <=  32'b00111110100010000010111111000101 ;
        3462:  q   <=  32'b00111110100010000011011101001101 ;
        3463:  q   <=  32'b00111110100010000011111011010101 ;
        3464:  q   <=  32'b00111110100010000100011001011101 ;
        3465:  q   <=  32'b00111110100010000100110111100101 ;
        3466:  q   <=  32'b00111110100010000101010101101100 ;
        3467:  q   <=  32'b00111110100010000101110011110011 ;
        3468:  q   <=  32'b00111110100010000110010001111001 ;
        3469:  q   <=  32'b00111110100010000110110000000000 ;
        3470:  q   <=  32'b00111110100010000111001110000110 ;
        3471:  q   <=  32'b00111110100010000111101100001100 ;
        3472:  q   <=  32'b00111110100010001000001010010010 ;
        3473:  q   <=  32'b00111110100010001000101000010111 ;
        3474:  q   <=  32'b00111110100010001001000110011100 ;
        3475:  q   <=  32'b00111110100010001001100100100001 ;
        3476:  q   <=  32'b00111110100010001010000010100110 ;
        3477:  q   <=  32'b00111110100010001010100000101010 ;
        3478:  q   <=  32'b00111110100010001010111110101110 ;
        3479:  q   <=  32'b00111110100010001011011100110010 ;
        3480:  q   <=  32'b00111110100010001011111010110110 ;
        3481:  q   <=  32'b00111110100010001100011000111001 ;
        3482:  q   <=  32'b00111110100010001100110110111100 ;
        3483:  q   <=  32'b00111110100010001101010100111111 ;
        3484:  q   <=  32'b00111110100010001101110011000010 ;
        3485:  q   <=  32'b00111110100010001110010001000100 ;
        3486:  q   <=  32'b00111110100010001110101111000110 ;
        3487:  q   <=  32'b00111110100010001111001101001000 ;
        3488:  q   <=  32'b00111110100010001111101011001010 ;
        3489:  q   <=  32'b00111110100010010000001001001011 ;
        3490:  q   <=  32'b00111110100010010000100111001100 ;
        3491:  q   <=  32'b00111110100010010001000101001101 ;
        3492:  q   <=  32'b00111110100010010001100011001110 ;
        3493:  q   <=  32'b00111110100010010010000001001110 ;
        3494:  q   <=  32'b00111110100010010010011111001110 ;
        3495:  q   <=  32'b00111110100010010010111101001110 ;
        3496:  q   <=  32'b00111110100010010011011011001101 ;
        3497:  q   <=  32'b00111110100010010011111001001101 ;
        3498:  q   <=  32'b00111110100010010100010111001100 ;
        3499:  q   <=  32'b00111110100010010100110101001011 ;
        3500:  q   <=  32'b00111110100010010101010011001001 ;
        3501:  q   <=  32'b00111110100010010101110001001000 ;
        3502:  q   <=  32'b00111110100010010110001111000110 ;
        3503:  q   <=  32'b00111110100010010110101101000011 ;
        3504:  q   <=  32'b00111110100010010111001011000001 ;
        3505:  q   <=  32'b00111110100010010111101000111110 ;
        3506:  q   <=  32'b00111110100010011000000110111011 ;
        3507:  q   <=  32'b00111110100010011000100100111000 ;
        3508:  q   <=  32'b00111110100010011001000010110101 ;
        3509:  q   <=  32'b00111110100010011001100000110001 ;
        3510:  q   <=  32'b00111110100010011001111110101101 ;
        3511:  q   <=  32'b00111110100010011010011100101001 ;
        3512:  q   <=  32'b00111110100010011010111010100100 ;
        3513:  q   <=  32'b00111110100010011011011000100000 ;
        3514:  q   <=  32'b00111110100010011011110110011011 ;
        3515:  q   <=  32'b00111110100010011100010100010110 ;
        3516:  q   <=  32'b00111110100010011100110010010000 ;
        3517:  q   <=  32'b00111110100010011101010000001010 ;
        3518:  q   <=  32'b00111110100010011101101110000100 ;
        3519:  q   <=  32'b00111110100010011110001011111110 ;
        3520:  q   <=  32'b00111110100010011110101001111000 ;
        3521:  q   <=  32'b00111110100010011111000111110001 ;
        3522:  q   <=  32'b00111110100010011111100101101010 ;
        3523:  q   <=  32'b00111110100010100000000011100011 ;
        3524:  q   <=  32'b00111110100010100000100001011011 ;
        3525:  q   <=  32'b00111110100010100000111111010100 ;
        3526:  q   <=  32'b00111110100010100001011101001100 ;
        3527:  q   <=  32'b00111110100010100001111011000011 ;
        3528:  q   <=  32'b00111110100010100010011000111011 ;
        3529:  q   <=  32'b00111110100010100010110110110010 ;
        3530:  q   <=  32'b00111110100010100011010100101001 ;
        3531:  q   <=  32'b00111110100010100011110010100000 ;
        3532:  q   <=  32'b00111110100010100100010000010111 ;
        3533:  q   <=  32'b00111110100010100100101110001101 ;
        3534:  q   <=  32'b00111110100010100101001100000011 ;
        3535:  q   <=  32'b00111110100010100101101001111001 ;
        3536:  q   <=  32'b00111110100010100110000111101110 ;
        3537:  q   <=  32'b00111110100010100110100101100011 ;
        3538:  q   <=  32'b00111110100010100111000011011000 ;
        3539:  q   <=  32'b00111110100010100111100001001101 ;
        3540:  q   <=  32'b00111110100010100111111111000010 ;
        3541:  q   <=  32'b00111110100010101000011100110110 ;
        3542:  q   <=  32'b00111110100010101000111010101010 ;
        3543:  q   <=  32'b00111110100010101001011000011110 ;
        3544:  q   <=  32'b00111110100010101001110110010001 ;
        3545:  q   <=  32'b00111110100010101010010100000101 ;
        3546:  q   <=  32'b00111110100010101010110001111000 ;
        3547:  q   <=  32'b00111110100010101011001111101010 ;
        3548:  q   <=  32'b00111110100010101011101101011101 ;
        3549:  q   <=  32'b00111110100010101100001011001111 ;
        3550:  q   <=  32'b00111110100010101100101001000001 ;
        3551:  q   <=  32'b00111110100010101101000110110011 ;
        3552:  q   <=  32'b00111110100010101101100100100101 ;
        3553:  q   <=  32'b00111110100010101110000010010110 ;
        3554:  q   <=  32'b00111110100010101110100000000111 ;
        3555:  q   <=  32'b00111110100010101110111101111000 ;
        3556:  q   <=  32'b00111110100010101111011011101000 ;
        3557:  q   <=  32'b00111110100010101111111001011000 ;
        3558:  q   <=  32'b00111110100010110000010111001000 ;
        3559:  q   <=  32'b00111110100010110000110100111000 ;
        3560:  q   <=  32'b00111110100010110001010010101000 ;
        3561:  q   <=  32'b00111110100010110001110000010111 ;
        3562:  q   <=  32'b00111110100010110010001110000110 ;
        3563:  q   <=  32'b00111110100010110010101011110101 ;
        3564:  q   <=  32'b00111110100010110011001001100011 ;
        3565:  q   <=  32'b00111110100010110011100111010010 ;
        3566:  q   <=  32'b00111110100010110100000101000000 ;
        3567:  q   <=  32'b00111110100010110100100010101110 ;
        3568:  q   <=  32'b00111110100010110101000000011011 ;
        3569:  q   <=  32'b00111110100010110101011110001000 ;
        3570:  q   <=  32'b00111110100010110101111011110101 ;
        3571:  q   <=  32'b00111110100010110110011001100010 ;
        3572:  q   <=  32'b00111110100010110110110111001111 ;
        3573:  q   <=  32'b00111110100010110111010100111011 ;
        3574:  q   <=  32'b00111110100010110111110010100111 ;
        3575:  q   <=  32'b00111110100010111000010000010011 ;
        3576:  q   <=  32'b00111110100010111000101101111111 ;
        3577:  q   <=  32'b00111110100010111001001011101010 ;
        3578:  q   <=  32'b00111110100010111001101001010101 ;
        3579:  q   <=  32'b00111110100010111010000111000000 ;
        3580:  q   <=  32'b00111110100010111010100100101010 ;
        3581:  q   <=  32'b00111110100010111011000010010101 ;
        3582:  q   <=  32'b00111110100010111011011111111111 ;
        3583:  q   <=  32'b00111110100010111011111101101001 ;
        3584:  q   <=  32'b00111110100010111100011011010010 ;
        3585:  q   <=  32'b00111110100010111100111000111011 ;
        3586:  q   <=  32'b00111110100010111101010110100101 ;
        3587:  q   <=  32'b00111110100010111101110100001101 ;
        3588:  q   <=  32'b00111110100010111110010001110110 ;
        3589:  q   <=  32'b00111110100010111110101111011110 ;
        3590:  q   <=  32'b00111110100010111111001101000110 ;
        3591:  q   <=  32'b00111110100010111111101010101110 ;
        3592:  q   <=  32'b00111110100011000000001000010110 ;
        3593:  q   <=  32'b00111110100011000000100101111101 ;
        3594:  q   <=  32'b00111110100011000001000011100100 ;
        3595:  q   <=  32'b00111110100011000001100001001011 ;
        3596:  q   <=  32'b00111110100011000001111110110010 ;
        3597:  q   <=  32'b00111110100011000010011100011000 ;
        3598:  q   <=  32'b00111110100011000010111001111110 ;
        3599:  q   <=  32'b00111110100011000011010111100100 ;
        3600:  q   <=  32'b00111110100011000011110101001010 ;
        3601:  q   <=  32'b00111110100011000100010010101111 ;
        3602:  q   <=  32'b00111110100011000100110000010100 ;
        3603:  q   <=  32'b00111110100011000101001101111001 ;
        3604:  q   <=  32'b00111110100011000101101011011110 ;
        3605:  q   <=  32'b00111110100011000110001001000010 ;
        3606:  q   <=  32'b00111110100011000110100110100111 ;
        3607:  q   <=  32'b00111110100011000111000100001011 ;
        3608:  q   <=  32'b00111110100011000111100001101110 ;
        3609:  q   <=  32'b00111110100011000111111111010010 ;
        3610:  q   <=  32'b00111110100011001000011100110101 ;
        3611:  q   <=  32'b00111110100011001000111010011000 ;
        3612:  q   <=  32'b00111110100011001001010111111010 ;
        3613:  q   <=  32'b00111110100011001001110101011101 ;
        3614:  q   <=  32'b00111110100011001010010010111111 ;
        3615:  q   <=  32'b00111110100011001010110000100001 ;
        3616:  q   <=  32'b00111110100011001011001110000011 ;
        3617:  q   <=  32'b00111110100011001011101011100100 ;
        3618:  q   <=  32'b00111110100011001100001001000101 ;
        3619:  q   <=  32'b00111110100011001100100110100110 ;
        3620:  q   <=  32'b00111110100011001101000100000111 ;
        3621:  q   <=  32'b00111110100011001101100001101000 ;
        3622:  q   <=  32'b00111110100011001101111111001000 ;
        3623:  q   <=  32'b00111110100011001110011100101000 ;
        3624:  q   <=  32'b00111110100011001110111010001000 ;
        3625:  q   <=  32'b00111110100011001111010111100111 ;
        3626:  q   <=  32'b00111110100011001111110101000110 ;
        3627:  q   <=  32'b00111110100011010000010010100101 ;
        3628:  q   <=  32'b00111110100011010000110000000100 ;
        3629:  q   <=  32'b00111110100011010001001101100011 ;
        3630:  q   <=  32'b00111110100011010001101011000001 ;
        3631:  q   <=  32'b00111110100011010010001000011111 ;
        3632:  q   <=  32'b00111110100011010010100101111101 ;
        3633:  q   <=  32'b00111110100011010011000011011010 ;
        3634:  q   <=  32'b00111110100011010011100000111000 ;
        3635:  q   <=  32'b00111110100011010011111110010101 ;
        3636:  q   <=  32'b00111110100011010100011011110010 ;
        3637:  q   <=  32'b00111110100011010100111001001110 ;
        3638:  q   <=  32'b00111110100011010101010110101011 ;
        3639:  q   <=  32'b00111110100011010101110100000111 ;
        3640:  q   <=  32'b00111110100011010110010001100010 ;
        3641:  q   <=  32'b00111110100011010110101110111110 ;
        3642:  q   <=  32'b00111110100011010111001100011001 ;
        3643:  q   <=  32'b00111110100011010111101001110101 ;
        3644:  q   <=  32'b00111110100011011000000111001111 ;
        3645:  q   <=  32'b00111110100011011000100100101010 ;
        3646:  q   <=  32'b00111110100011011001000010000100 ;
        3647:  q   <=  32'b00111110100011011001011111011111 ;
        3648:  q   <=  32'b00111110100011011001111100111000 ;
        3649:  q   <=  32'b00111110100011011010011010010010 ;
        3650:  q   <=  32'b00111110100011011010110111101100 ;
        3651:  q   <=  32'b00111110100011011011010101000101 ;
        3652:  q   <=  32'b00111110100011011011110010011110 ;
        3653:  q   <=  32'b00111110100011011100001111110110 ;
        3654:  q   <=  32'b00111110100011011100101101001111 ;
        3655:  q   <=  32'b00111110100011011101001010100111 ;
        3656:  q   <=  32'b00111110100011011101100111111111 ;
        3657:  q   <=  32'b00111110100011011110000101010111 ;
        3658:  q   <=  32'b00111110100011011110100010101110 ;
        3659:  q   <=  32'b00111110100011011111000000000101 ;
        3660:  q   <=  32'b00111110100011011111011101011100 ;
        3661:  q   <=  32'b00111110100011011111111010110011 ;
        3662:  q   <=  32'b00111110100011100000011000001010 ;
        3663:  q   <=  32'b00111110100011100000110101100000 ;
        3664:  q   <=  32'b00111110100011100001010010110110 ;
        3665:  q   <=  32'b00111110100011100001110000001100 ;
        3666:  q   <=  32'b00111110100011100010001101100001 ;
        3667:  q   <=  32'b00111110100011100010101010110110 ;
        3668:  q   <=  32'b00111110100011100011001000001100 ;
        3669:  q   <=  32'b00111110100011100011100101100000 ;
        3670:  q   <=  32'b00111110100011100100000010110101 ;
        3671:  q   <=  32'b00111110100011100100100000001001 ;
        3672:  q   <=  32'b00111110100011100100111101011101 ;
        3673:  q   <=  32'b00111110100011100101011010110001 ;
        3674:  q   <=  32'b00111110100011100101111000000101 ;
        3675:  q   <=  32'b00111110100011100110010101011000 ;
        3676:  q   <=  32'b00111110100011100110110010101011 ;
        3677:  q   <=  32'b00111110100011100111001111111110 ;
        3678:  q   <=  32'b00111110100011100111101101010001 ;
        3679:  q   <=  32'b00111110100011101000001010100011 ;
        3680:  q   <=  32'b00111110100011101000100111110101 ;
        3681:  q   <=  32'b00111110100011101001000101000111 ;
        3682:  q   <=  32'b00111110100011101001100010011001 ;
        3683:  q   <=  32'b00111110100011101001111111101010 ;
        3684:  q   <=  32'b00111110100011101010011100111100 ;
        3685:  q   <=  32'b00111110100011101010111010001101 ;
        3686:  q   <=  32'b00111110100011101011010111011101 ;
        3687:  q   <=  32'b00111110100011101011110100101110 ;
        3688:  q   <=  32'b00111110100011101100010001111110 ;
        3689:  q   <=  32'b00111110100011101100101111001110 ;
        3690:  q   <=  32'b00111110100011101101001100011110 ;
        3691:  q   <=  32'b00111110100011101101101001101101 ;
        3692:  q   <=  32'b00111110100011101110000110111100 ;
        3693:  q   <=  32'b00111110100011101110100100001011 ;
        3694:  q   <=  32'b00111110100011101111000001011010 ;
        3695:  q   <=  32'b00111110100011101111011110101001 ;
        3696:  q   <=  32'b00111110100011101111111011110111 ;
        3697:  q   <=  32'b00111110100011110000011001000101 ;
        3698:  q   <=  32'b00111110100011110000110110010011 ;
        3699:  q   <=  32'b00111110100011110001010011100001 ;
        3700:  q   <=  32'b00111110100011110001110000101110 ;
        3701:  q   <=  32'b00111110100011110010001101111011 ;
        3702:  q   <=  32'b00111110100011110010101011001000 ;
        3703:  q   <=  32'b00111110100011110011001000010101 ;
        3704:  q   <=  32'b00111110100011110011100101100001 ;
        3705:  q   <=  32'b00111110100011110100000010101101 ;
        3706:  q   <=  32'b00111110100011110100011111111001 ;
        3707:  q   <=  32'b00111110100011110100111101000101 ;
        3708:  q   <=  32'b00111110100011110101011010010000 ;
        3709:  q   <=  32'b00111110100011110101110111011011 ;
        3710:  q   <=  32'b00111110100011110110010100100110 ;
        3711:  q   <=  32'b00111110100011110110110001110001 ;
        3712:  q   <=  32'b00111110100011110111001110111011 ;
        3713:  q   <=  32'b00111110100011110111101100000110 ;
        3714:  q   <=  32'b00111110100011111000001001010000 ;
        3715:  q   <=  32'b00111110100011111000100110011001 ;
        3716:  q   <=  32'b00111110100011111001000011100011 ;
        3717:  q   <=  32'b00111110100011111001100000101100 ;
        3718:  q   <=  32'b00111110100011111001111101110101 ;
        3719:  q   <=  32'b00111110100011111010011010111110 ;
        3720:  q   <=  32'b00111110100011111010111000000111 ;
        3721:  q   <=  32'b00111110100011111011010101001111 ;
        3722:  q   <=  32'b00111110100011111011110010010111 ;
        3723:  q   <=  32'b00111110100011111100001111011111 ;
        3724:  q   <=  32'b00111110100011111100101100100111 ;
        3725:  q   <=  32'b00111110100011111101001001101110 ;
        3726:  q   <=  32'b00111110100011111101100110110101 ;
        3727:  q   <=  32'b00111110100011111110000011111100 ;
        3728:  q   <=  32'b00111110100011111110100001000011 ;
        3729:  q   <=  32'b00111110100011111110111110001001 ;
        3730:  q   <=  32'b00111110100011111111011011001111 ;
        3731:  q   <=  32'b00111110100011111111111000010101 ;
        3732:  q   <=  32'b00111110100100000000010101011011 ;
        3733:  q   <=  32'b00111110100100000000110010100000 ;
        3734:  q   <=  32'b00111110100100000001001111100110 ;
        3735:  q   <=  32'b00111110100100000001101100101011 ;
        3736:  q   <=  32'b00111110100100000010001001101111 ;
        3737:  q   <=  32'b00111110100100000010100110110100 ;
        3738:  q   <=  32'b00111110100100000011000011111000 ;
        3739:  q   <=  32'b00111110100100000011100000111100 ;
        3740:  q   <=  32'b00111110100100000011111110000000 ;
        3741:  q   <=  32'b00111110100100000100011011000011 ;
        3742:  q   <=  32'b00111110100100000100111000000111 ;
        3743:  q   <=  32'b00111110100100000101010101001010 ;
        3744:  q   <=  32'b00111110100100000101110010001101 ;
        3745:  q   <=  32'b00111110100100000110001111001111 ;
        3746:  q   <=  32'b00111110100100000110101100010010 ;
        3747:  q   <=  32'b00111110100100000111001001010100 ;
        3748:  q   <=  32'b00111110100100000111100110010110 ;
        3749:  q   <=  32'b00111110100100001000000011011000 ;
        3750:  q   <=  32'b00111110100100001000100000011001 ;
        3751:  q   <=  32'b00111110100100001000111101011010 ;
        3752:  q   <=  32'b00111110100100001001011010011011 ;
        3753:  q   <=  32'b00111110100100001001110111011100 ;
        3754:  q   <=  32'b00111110100100001010010100011100 ;
        3755:  q   <=  32'b00111110100100001010110001011101 ;
        3756:  q   <=  32'b00111110100100001011001110011101 ;
        3757:  q   <=  32'b00111110100100001011101011011100 ;
        3758:  q   <=  32'b00111110100100001100001000011100 ;
        3759:  q   <=  32'b00111110100100001100100101011011 ;
        3760:  q   <=  32'b00111110100100001101000010011010 ;
        3761:  q   <=  32'b00111110100100001101011111011001 ;
        3762:  q   <=  32'b00111110100100001101111100011000 ;
        3763:  q   <=  32'b00111110100100001110011001010110 ;
        3764:  q   <=  32'b00111110100100001110110110010100 ;
        3765:  q   <=  32'b00111110100100001111010011010010 ;
        3766:  q   <=  32'b00111110100100001111110000010000 ;
        3767:  q   <=  32'b00111110100100010000001101001101 ;
        3768:  q   <=  32'b00111110100100010000101010001010 ;
        3769:  q   <=  32'b00111110100100010001000111000111 ;
        3770:  q   <=  32'b00111110100100010001100100000100 ;
        3771:  q   <=  32'b00111110100100010010000001000000 ;
        3772:  q   <=  32'b00111110100100010010011101111101 ;
        3773:  q   <=  32'b00111110100100010010111010111001 ;
        3774:  q   <=  32'b00111110100100010011010111110100 ;
        3775:  q   <=  32'b00111110100100010011110100110000 ;
        3776:  q   <=  32'b00111110100100010100010001101011 ;
        3777:  q   <=  32'b00111110100100010100101110100110 ;
        3778:  q   <=  32'b00111110100100010101001011100001 ;
        3779:  q   <=  32'b00111110100100010101101000011100 ;
        3780:  q   <=  32'b00111110100100010110000101010110 ;
        3781:  q   <=  32'b00111110100100010110100010010000 ;
        3782:  q   <=  32'b00111110100100010110111111001010 ;
        3783:  q   <=  32'b00111110100100010111011100000100 ;
        3784:  q   <=  32'b00111110100100010111111000111101 ;
        3785:  q   <=  32'b00111110100100011000010101110110 ;
        3786:  q   <=  32'b00111110100100011000110010101111 ;
        3787:  q   <=  32'b00111110100100011001001111101000 ;
        3788:  q   <=  32'b00111110100100011001101100100001 ;
        3789:  q   <=  32'b00111110100100011010001001011001 ;
        3790:  q   <=  32'b00111110100100011010100110010001 ;
        3791:  q   <=  32'b00111110100100011011000011001001 ;
        3792:  q   <=  32'b00111110100100011011100000000000 ;
        3793:  q   <=  32'b00111110100100011011111100110111 ;
        3794:  q   <=  32'b00111110100100011100011001101111 ;
        3795:  q   <=  32'b00111110100100011100110110100101 ;
        3796:  q   <=  32'b00111110100100011101010011011100 ;
        3797:  q   <=  32'b00111110100100011101110000010010 ;
        3798:  q   <=  32'b00111110100100011110001101001001 ;
        3799:  q   <=  32'b00111110100100011110101001111110 ;
        3800:  q   <=  32'b00111110100100011111000110110100 ;
        3801:  q   <=  32'b00111110100100011111100011101010 ;
        3802:  q   <=  32'b00111110100100100000000000011111 ;
        3803:  q   <=  32'b00111110100100100000011101010100 ;
        3804:  q   <=  32'b00111110100100100000111010001000 ;
        3805:  q   <=  32'b00111110100100100001010110111101 ;
        3806:  q   <=  32'b00111110100100100001110011110001 ;
        3807:  q   <=  32'b00111110100100100010010000100101 ;
        3808:  q   <=  32'b00111110100100100010101101011001 ;
        3809:  q   <=  32'b00111110100100100011001010001101 ;
        3810:  q   <=  32'b00111110100100100011100111000000 ;
        3811:  q   <=  32'b00111110100100100100000011110011 ;
        3812:  q   <=  32'b00111110100100100100100000100110 ;
        3813:  q   <=  32'b00111110100100100100111101011001 ;
        3814:  q   <=  32'b00111110100100100101011010001011 ;
        3815:  q   <=  32'b00111110100100100101110110111101 ;
        3816:  q   <=  32'b00111110100100100110010011101111 ;
        3817:  q   <=  32'b00111110100100100110110000100001 ;
        3818:  q   <=  32'b00111110100100100111001101010010 ;
        3819:  q   <=  32'b00111110100100100111101010000100 ;
        3820:  q   <=  32'b00111110100100101000000110110101 ;
        3821:  q   <=  32'b00111110100100101000100011100101 ;
        3822:  q   <=  32'b00111110100100101001000000010110 ;
        3823:  q   <=  32'b00111110100100101001011101000110 ;
        3824:  q   <=  32'b00111110100100101001111001110110 ;
        3825:  q   <=  32'b00111110100100101010010110100110 ;
        3826:  q   <=  32'b00111110100100101010110011010110 ;
        3827:  q   <=  32'b00111110100100101011010000000101 ;
        3828:  q   <=  32'b00111110100100101011101100110100 ;
        3829:  q   <=  32'b00111110100100101100001001100011 ;
        3830:  q   <=  32'b00111110100100101100100110010010 ;
        3831:  q   <=  32'b00111110100100101101000011000000 ;
        3832:  q   <=  32'b00111110100100101101011111101111 ;
        3833:  q   <=  32'b00111110100100101101111100011101 ;
        3834:  q   <=  32'b00111110100100101110011001001010 ;
        3835:  q   <=  32'b00111110100100101110110101111000 ;
        3836:  q   <=  32'b00111110100100101111010010100101 ;
        3837:  q   <=  32'b00111110100100101111101111010010 ;
        3838:  q   <=  32'b00111110100100110000001011111111 ;
        3839:  q   <=  32'b00111110100100110000101000101100 ;
        3840:  q   <=  32'b00111110100100110001000101011000 ;
        3841:  q   <=  32'b00111110100100110001100010000100 ;
        3842:  q   <=  32'b00111110100100110001111110110000 ;
        3843:  q   <=  32'b00111110100100110010011011011100 ;
        3844:  q   <=  32'b00111110100100110010111000000111 ;
        3845:  q   <=  32'b00111110100100110011010100110010 ;
        3846:  q   <=  32'b00111110100100110011110001011101 ;
        3847:  q   <=  32'b00111110100100110100001110001000 ;
        3848:  q   <=  32'b00111110100100110100101010110011 ;
        3849:  q   <=  32'b00111110100100110101000111011101 ;
        3850:  q   <=  32'b00111110100100110101100100000111 ;
        3851:  q   <=  32'b00111110100100110110000000110001 ;
        3852:  q   <=  32'b00111110100100110110011101011010 ;
        3853:  q   <=  32'b00111110100100110110111010000100 ;
        3854:  q   <=  32'b00111110100100110111010110101101 ;
        3855:  q   <=  32'b00111110100100110111110011010110 ;
        3856:  q   <=  32'b00111110100100111000001111111110 ;
        3857:  q   <=  32'b00111110100100111000101100100111 ;
        3858:  q   <=  32'b00111110100100111001001001001111 ;
        3859:  q   <=  32'b00111110100100111001100101110111 ;
        3860:  q   <=  32'b00111110100100111010000010011111 ;
        3861:  q   <=  32'b00111110100100111010011111000110 ;
        3862:  q   <=  32'b00111110100100111010111011101110 ;
        3863:  q   <=  32'b00111110100100111011011000010101 ;
        3864:  q   <=  32'b00111110100100111011110100111100 ;
        3865:  q   <=  32'b00111110100100111100010001100010 ;
        3866:  q   <=  32'b00111110100100111100101110001001 ;
        3867:  q   <=  32'b00111110100100111101001010101111 ;
        3868:  q   <=  32'b00111110100100111101100111010101 ;
        3869:  q   <=  32'b00111110100100111110000011111010 ;
        3870:  q   <=  32'b00111110100100111110100000100000 ;
        3871:  q   <=  32'b00111110100100111110111101000101 ;
        3872:  q   <=  32'b00111110100100111111011001101010 ;
        3873:  q   <=  32'b00111110100100111111110110001111 ;
        3874:  q   <=  32'b00111110100101000000010010110011 ;
        3875:  q   <=  32'b00111110100101000000101111011000 ;
        3876:  q   <=  32'b00111110100101000001001011111100 ;
        3877:  q   <=  32'b00111110100101000001101000011111 ;
        3878:  q   <=  32'b00111110100101000010000101000011 ;
        3879:  q   <=  32'b00111110100101000010100001100110 ;
        3880:  q   <=  32'b00111110100101000010111110001010 ;
        3881:  q   <=  32'b00111110100101000011011010101101 ;
        3882:  q   <=  32'b00111110100101000011110111001111 ;
        3883:  q   <=  32'b00111110100101000100010011110010 ;
        3884:  q   <=  32'b00111110100101000100110000010100 ;
        3885:  q   <=  32'b00111110100101000101001100110110 ;
        3886:  q   <=  32'b00111110100101000101101001011000 ;
        3887:  q   <=  32'b00111110100101000110000101111001 ;
        3888:  q   <=  32'b00111110100101000110100010011011 ;
        3889:  q   <=  32'b00111110100101000110111110111100 ;
        3890:  q   <=  32'b00111110100101000111011011011101 ;
        3891:  q   <=  32'b00111110100101000111110111111101 ;
        3892:  q   <=  32'b00111110100101001000010100011110 ;
        3893:  q   <=  32'b00111110100101001000110000111110 ;
        3894:  q   <=  32'b00111110100101001001001101011110 ;
        3895:  q   <=  32'b00111110100101001001101001111110 ;
        3896:  q   <=  32'b00111110100101001010000110011101 ;
        3897:  q   <=  32'b00111110100101001010100010111100 ;
        3898:  q   <=  32'b00111110100101001010111111011011 ;
        3899:  q   <=  32'b00111110100101001011011011111010 ;
        3900:  q   <=  32'b00111110100101001011111000011001 ;
        3901:  q   <=  32'b00111110100101001100010100110111 ;
        3902:  q   <=  32'b00111110100101001100110001010101 ;
        3903:  q   <=  32'b00111110100101001101001101110011 ;
        3904:  q   <=  32'b00111110100101001101101010010001 ;
        3905:  q   <=  32'b00111110100101001110000110101110 ;
        3906:  q   <=  32'b00111110100101001110100011001011 ;
        3907:  q   <=  32'b00111110100101001110111111101000 ;
        3908:  q   <=  32'b00111110100101001111011100000101 ;
        3909:  q   <=  32'b00111110100101001111111000100010 ;
        3910:  q   <=  32'b00111110100101010000010100111110 ;
        3911:  q   <=  32'b00111110100101010000110001011010 ;
        3912:  q   <=  32'b00111110100101010001001101110110 ;
        3913:  q   <=  32'b00111110100101010001101010010010 ;
        3914:  q   <=  32'b00111110100101010010000110101101 ;
        3915:  q   <=  32'b00111110100101010010100011001000 ;
        3916:  q   <=  32'b00111110100101010010111111100011 ;
        3917:  q   <=  32'b00111110100101010011011011111110 ;
        3918:  q   <=  32'b00111110100101010011111000011000 ;
        3919:  q   <=  32'b00111110100101010100010100110011 ;
        3920:  q   <=  32'b00111110100101010100110001001101 ;
        3921:  q   <=  32'b00111110100101010101001101100111 ;
        3922:  q   <=  32'b00111110100101010101101010000000 ;
        3923:  q   <=  32'b00111110100101010110000110011001 ;
        3924:  q   <=  32'b00111110100101010110100010110011 ;
        3925:  q   <=  32'b00111110100101010110111111001100 ;
        3926:  q   <=  32'b00111110100101010111011011100100 ;
        3927:  q   <=  32'b00111110100101010111110111111101 ;
        3928:  q   <=  32'b00111110100101011000010100010101 ;
        3929:  q   <=  32'b00111110100101011000110000101101 ;
        3930:  q   <=  32'b00111110100101011001001101000101 ;
        3931:  q   <=  32'b00111110100101011001101001011100 ;
        3932:  q   <=  32'b00111110100101011010000101110100 ;
        3933:  q   <=  32'b00111110100101011010100010001011 ;
        3934:  q   <=  32'b00111110100101011010111110100010 ;
        3935:  q   <=  32'b00111110100101011011011010111000 ;
        3936:  q   <=  32'b00111110100101011011110111001111 ;
        3937:  q   <=  32'b00111110100101011100010011100101 ;
        3938:  q   <=  32'b00111110100101011100101111111011 ;
        3939:  q   <=  32'b00111110100101011101001100010000 ;
        3940:  q   <=  32'b00111110100101011101101000100110 ;
        3941:  q   <=  32'b00111110100101011110000100111011 ;
        3942:  q   <=  32'b00111110100101011110100001010000 ;
        3943:  q   <=  32'b00111110100101011110111101100101 ;
        3944:  q   <=  32'b00111110100101011111011001111010 ;
        3945:  q   <=  32'b00111110100101011111110110001110 ;
        3946:  q   <=  32'b00111110100101100000010010100010 ;
        3947:  q   <=  32'b00111110100101100000101110110110 ;
        3948:  q   <=  32'b00111110100101100001001011001010 ;
        3949:  q   <=  32'b00111110100101100001100111011101 ;
        3950:  q   <=  32'b00111110100101100010000011110001 ;
        3951:  q   <=  32'b00111110100101100010100000000100 ;
        3952:  q   <=  32'b00111110100101100010111100010111 ;
        3953:  q   <=  32'b00111110100101100011011000101001 ;
        3954:  q   <=  32'b00111110100101100011110100111100 ;
        3955:  q   <=  32'b00111110100101100100010001001110 ;
        3956:  q   <=  32'b00111110100101100100101101100000 ;
        3957:  q   <=  32'b00111110100101100101001001110001 ;
        3958:  q   <=  32'b00111110100101100101100110000011 ;
        3959:  q   <=  32'b00111110100101100110000010010100 ;
        3960:  q   <=  32'b00111110100101100110011110100101 ;
        3961:  q   <=  32'b00111110100101100110111010110110 ;
        3962:  q   <=  32'b00111110100101100111010111000110 ;
        3963:  q   <=  32'b00111110100101100111110011010111 ;
        3964:  q   <=  32'b00111110100101101000001111100111 ;
        3965:  q   <=  32'b00111110100101101000101011110111 ;
        3966:  q   <=  32'b00111110100101101001001000000110 ;
        3967:  q   <=  32'b00111110100101101001100100010110 ;
        3968:  q   <=  32'b00111110100101101010000000100101 ;
        3969:  q   <=  32'b00111110100101101010011100110100 ;
        3970:  q   <=  32'b00111110100101101010111001000011 ;
        3971:  q   <=  32'b00111110100101101011010101010001 ;
        3972:  q   <=  32'b00111110100101101011110001100000 ;
        3973:  q   <=  32'b00111110100101101100001101101110 ;
        3974:  q   <=  32'b00111110100101101100101001111100 ;
        3975:  q   <=  32'b00111110100101101101000110001001 ;
        3976:  q   <=  32'b00111110100101101101100010010111 ;
        3977:  q   <=  32'b00111110100101101101111110100100 ;
        3978:  q   <=  32'b00111110100101101110011010110001 ;
        3979:  q   <=  32'b00111110100101101110110110111110 ;
        3980:  q   <=  32'b00111110100101101111010011001010 ;
        3981:  q   <=  32'b00111110100101101111101111010110 ;
        3982:  q   <=  32'b00111110100101110000001011100011 ;
        3983:  q   <=  32'b00111110100101110000100111101110 ;
        3984:  q   <=  32'b00111110100101110001000011111010 ;
        3985:  q   <=  32'b00111110100101110001100000000101 ;
        3986:  q   <=  32'b00111110100101110001111100010001 ;
        3987:  q   <=  32'b00111110100101110010011000011100 ;
        3988:  q   <=  32'b00111110100101110010110100100110 ;
        3989:  q   <=  32'b00111110100101110011010000110001 ;
        3990:  q   <=  32'b00111110100101110011101100111011 ;
        3991:  q   <=  32'b00111110100101110100001001000101 ;
        3992:  q   <=  32'b00111110100101110100100101001111 ;
        3993:  q   <=  32'b00111110100101110101000001011001 ;
        3994:  q   <=  32'b00111110100101110101011101100010 ;
        3995:  q   <=  32'b00111110100101110101111001101011 ;
        3996:  q   <=  32'b00111110100101110110010101110100 ;
        3997:  q   <=  32'b00111110100101110110110001111101 ;
        3998:  q   <=  32'b00111110100101110111001110000110 ;
        3999:  q   <=  32'b00111110100101110111101010001110 ;
        4000:  q   <=  32'b00111110100101111000000110010110 ;
        4001:  q   <=  32'b00111110100101111000100010011110 ;
        4002:  q   <=  32'b00111110100101111000111110100101 ;
        4003:  q   <=  32'b00111110100101111001011010101101 ;
        4004:  q   <=  32'b00111110100101111001110110110100 ;
        4005:  q   <=  32'b00111110100101111010010010111011 ;
        4006:  q   <=  32'b00111110100101111010101111000010 ;
        4007:  q   <=  32'b00111110100101111011001011001000 ;
        4008:  q   <=  32'b00111110100101111011100111001111 ;
        4009:  q   <=  32'b00111110100101111100000011010101 ;
        4010:  q   <=  32'b00111110100101111100011111011011 ;
        4011:  q   <=  32'b00111110100101111100111011100000 ;
        4012:  q   <=  32'b00111110100101111101010111100110 ;
        4013:  q   <=  32'b00111110100101111101110011101011 ;
        4014:  q   <=  32'b00111110100101111110001111110000 ;
        4015:  q   <=  32'b00111110100101111110101011110100 ;
        4016:  q   <=  32'b00111110100101111111000111111001 ;
        4017:  q   <=  32'b00111110100101111111100011111101 ;
        4018:  q   <=  32'b00111110100110000000000000000001 ;
        4019:  q   <=  32'b00111110100110000000011100000101 ;
        4020:  q   <=  32'b00111110100110000000111000001001 ;
        4021:  q   <=  32'b00111110100110000001010100001100 ;
        4022:  q   <=  32'b00111110100110000001110000001111 ;
        4023:  q   <=  32'b00111110100110000010001100010010 ;
        4024:  q   <=  32'b00111110100110000010101000010101 ;
        4025:  q   <=  32'b00111110100110000011000100011000 ;
        4026:  q   <=  32'b00111110100110000011100000011010 ;
        4027:  q   <=  32'b00111110100110000011111100011100 ;
        4028:  q   <=  32'b00111110100110000100011000011110 ;
        4029:  q   <=  32'b00111110100110000100110100100000 ;
        4030:  q   <=  32'b00111110100110000101010000100001 ;
        4031:  q   <=  32'b00111110100110000101101100100010 ;
        4032:  q   <=  32'b00111110100110000110001000100011 ;
        4033:  q   <=  32'b00111110100110000110100100100100 ;
        4034:  q   <=  32'b00111110100110000111000000100101 ;
        4035:  q   <=  32'b00111110100110000111011100100101 ;
        4036:  q   <=  32'b00111110100110000111111000100101 ;
        4037:  q   <=  32'b00111110100110001000010100100101 ;
        4038:  q   <=  32'b00111110100110001000110000100101 ;
        4039:  q   <=  32'b00111110100110001001001100100100 ;
        4040:  q   <=  32'b00111110100110001001101000100011 ;
        4041:  q   <=  32'b00111110100110001010000100100010 ;
        4042:  q   <=  32'b00111110100110001010100000100001 ;
        4043:  q   <=  32'b00111110100110001010111100100000 ;
        4044:  q   <=  32'b00111110100110001011011000011110 ;
        4045:  q   <=  32'b00111110100110001011110100011100 ;
        4046:  q   <=  32'b00111110100110001100010000011010 ;
        4047:  q   <=  32'b00111110100110001100101100011000 ;
        4048:  q   <=  32'b00111110100110001101001000010101 ;
        4049:  q   <=  32'b00111110100110001101100100010010 ;
        4050:  q   <=  32'b00111110100110001110000000001111 ;
        4051:  q   <=  32'b00111110100110001110011100001100 ;
        4052:  q   <=  32'b00111110100110001110111000001001 ;
        4053:  q   <=  32'b00111110100110001111010100000101 ;
        4054:  q   <=  32'b00111110100110001111110000000001 ;
        4055:  q   <=  32'b00111110100110010000001011111101 ;
        4056:  q   <=  32'b00111110100110010000100111111001 ;
        4057:  q   <=  32'b00111110100110010001000011110100 ;
        4058:  q   <=  32'b00111110100110010001011111110000 ;
        4059:  q   <=  32'b00111110100110010001111011101011 ;
        4060:  q   <=  32'b00111110100110010010010111100110 ;
        4061:  q   <=  32'b00111110100110010010110011100000 ;
        4062:  q   <=  32'b00111110100110010011001111011011 ;
        4063:  q   <=  32'b00111110100110010011101011010101 ;
        4064:  q   <=  32'b00111110100110010100000111001111 ;
        4065:  q   <=  32'b00111110100110010100100011001000 ;
        4066:  q   <=  32'b00111110100110010100111111000010 ;
        4067:  q   <=  32'b00111110100110010101011010111011 ;
        4068:  q   <=  32'b00111110100110010101110110110100 ;
        4069:  q   <=  32'b00111110100110010110010010101101 ;
        4070:  q   <=  32'b00111110100110010110101110100110 ;
        4071:  q   <=  32'b00111110100110010111001010011110 ;
        4072:  q   <=  32'b00111110100110010111100110010110 ;
        4073:  q   <=  32'b00111110100110011000000010001110 ;
        4074:  q   <=  32'b00111110100110011000011110000110 ;
        4075:  q   <=  32'b00111110100110011000111001111110 ;
        4076:  q   <=  32'b00111110100110011001010101110101 ;
        4077:  q   <=  32'b00111110100110011001110001101100 ;
        4078:  q   <=  32'b00111110100110011010001101100011 ;
        4079:  q   <=  32'b00111110100110011010101001011010 ;
        4080:  q   <=  32'b00111110100110011011000101010000 ;
        4081:  q   <=  32'b00111110100110011011100001000111 ;
        4082:  q   <=  32'b00111110100110011011111100111101 ;
        4083:  q   <=  32'b00111110100110011100011000110010 ;
        4084:  q   <=  32'b00111110100110011100110100101000 ;
        4085:  q   <=  32'b00111110100110011101010000011101 ;
        4086:  q   <=  32'b00111110100110011101101100010010 ;
        4087:  q   <=  32'b00111110100110011110001000000111 ;
        4088:  q   <=  32'b00111110100110011110100011111100 ;
        4089:  q   <=  32'b00111110100110011110111111110001 ;
        4090:  q   <=  32'b00111110100110011111011011100101 ;
        4091:  q   <=  32'b00111110100110011111110111011001 ;
        4092:  q   <=  32'b00111110100110100000010011001101 ;
        4093:  q   <=  32'b00111110100110100000101111000000 ;
        4094:  q   <=  32'b00111110100110100001001010110100 ;
        4095:  q   <=  32'b00111110100110100001100110100111;
        default: q <= 0;
    endcase
end
endmodule
