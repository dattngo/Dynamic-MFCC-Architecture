module mem_w_image (clk, addr, cen, wen, data,q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00000000000000000000000000000000 ;
        2:  q   <=  32'b10111100010010010000111010001111 ;
        3:  q   <=  32'b10111100110010010000101010101111 ;
        4:  q   <=  32'b10111101000101101100001100101011 ;
        5:  q   <=  32'b10111101010010001111101100101111 ;
        6:  q   <=  32'b10111101011110110010101101110011 ;
        7:  q   <=  32'b10111101100101101010100100000100 ;
        8:  q   <=  32'b10111101101011111011011010000000 ;
        9:  q   <=  32'b10111101110010001011110100110101 ;
        10:  q   <=  32'b10111101111000011011110000101110 ;
        11:  q   <=  32'b10111101111110101011001001110010 ;
        12:  q   <=  32'b10111110000010011100111110000110 ;
        13:  q   <=  32'b10111110000101100100000010000011 ;
        14:  q   <=  32'b10111110001000101010101110110101 ;
        15:  q   <=  32'b10111110001011110001000010100010 ;
        16:  q   <=  32'b10111110001110110110111011001110 ;
        17:  q   <=  32'b10111110010001111100010111000001 ;
        18:  q   <=  32'b10111110010101000001010100000001 ;
        19:  q   <=  32'b10111110011000000101110000010011 ;
        20:  q   <=  32'b10111110011011001001101001111111 ;
        21:  q   <=  32'b10111110011110001100111111001011 ;
        22:  q   <=  32'b10111110100000100111110111000000 ;
        23:  q   <=  32'b10111110100010001000111010010011 ;
        24:  q   <=  32'b10111110100011101001101000100001 ;
        25:  q   <=  32'b10111110100101001010000000110001 ;
        26:  q   <=  32'b10111110100110101010000010000110 ;
        27:  q   <=  32'b10111110101000001001101011100100 ;
        28:  q   <=  32'b10111110101001101000111100010010 ;
        29:  q   <=  32'b10111110101011000111110011010011 ;
        30:  q   <=  32'b10111110101100100110001111101110 ;
        31:  q   <=  32'b10111110101110000100010000101001 ;
        32:  q   <=  32'b10111110101111100001110101001001 ;
        33:  q   <=  32'b10111110110000111110111100010101 ;
        34:  q   <=  32'b10111110110010011011100101010011 ;
        35:  q   <=  32'b10111110110011110111101111001010 ;
        36:  q   <=  32'b10111110110101010011011001000001 ;
        37:  q   <=  32'b10111110110110101110100010000000 ;
        38:  q   <=  32'b10111110111000001001001001001110 ;
        39:  q   <=  32'b10111110111001100011001101110100 ;
        40:  q   <=  32'b10111110111010111100101110111010 ;
        41:  q   <=  32'b10111110111100010101101011101001 ;
        42:  q   <=  32'b10111110111101101110000011001010 ;
        43:  q   <=  32'b10111110111111000101110100100110 ;
        44:  q   <=  32'b10111111000000001110011111100100 ;
        45:  q   <=  32'b10111111000000111001110000111100 ;
        46:  q   <=  32'b10111111000001100100101110000010 ;
        47:  q   <=  32'b10111111000010001111010110011010 ;
        48:  q   <=  32'b10111111000010111001101001101011 ;
        49:  q   <=  32'b10111111000011100011100111011001 ;
        50:  q   <=  32'b10111111000100001101001111001100 ;
        51:  q   <=  32'b10111111000100110110100000101010 ;
        52:  q   <=  32'b10111111000101011111011011011001 ;
        53:  q   <=  32'b10111111000110000111111110111111 ;
        54:  q   <=  32'b10111111000110110000001011000101 ;
        55:  q   <=  32'b10111111000111010111111111010001 ;
        56:  q   <=  32'b10111111000111111111011011001010 ;
        57:  q   <=  32'b10111111001000100110011110011001 ;
        58:  q   <=  32'b10111111001001001101001000100100 ;
        59:  q   <=  32'b10111111001001110011011001010101 ;
        60:  q   <=  32'b10111111001010011001010000010100 ;
        61:  q   <=  32'b10111111001010111110101101001001 ;
        62:  q   <=  32'b10111111001011100011101111011101 ;
        63:  q   <=  32'b10111111001100001000010110111010 ;
        64:  q   <=  32'b10111111001100101100100011001001 ;
        65:  q   <=  32'b10111111001101010000010011110011 ;
        66:  q   <=  32'b10111111001101110011101000100010 ;
        67:  q   <=  32'b10111111001110010110100001000001 ;
        68:  q   <=  32'b10111111001110111000111100111010 ;
        69:  q   <=  32'b10111111001111011010111011111001 ;
        70:  q   <=  32'b10111111001111111100011101100111 ;
        71:  q   <=  32'b10111111010000011101100001110000 ;
        72:  q   <=  32'b10111111010000111110001000000000 ;
        73:  q   <=  32'b10111111010001011110010000000011 ;
        74:  q   <=  32'b10111111010001111101111001100101 ;
        75:  q   <=  32'b10111111010010011101000100010010 ;
        76:  q   <=  32'b10111111010010111011101111110111 ;
        77:  q   <=  32'b10111111010011011001111100000010 ;
        78:  q   <=  32'b10111111010011110111101000011111 ;
        79:  q   <=  32'b10111111010100010100110100111101 ;
        80:  q   <=  32'b10111111010100110001100001001000 ;
        81:  q   <=  32'b10111111010101001101101100110001 ;
        82:  q   <=  32'b10111111010101101001010111100100 ;
        83:  q   <=  32'b10111111010110000100100001010010 ;
        84:  q   <=  32'b10111111010110011111001001101001 ;
        85:  q   <=  32'b10111111010110111001010000011010 ;
        86:  q   <=  32'b10111111010111010010110101010011 ;
        87:  q   <=  32'b10111111010111101011111000000101 ;
        88:  q   <=  32'b10111111011000000100011000100001 ;
        89:  q   <=  32'b10111111011000011100010110010111 ;
        90:  q   <=  32'b10111111011000110011110001011001 ;
        91:  q   <=  32'b10111111011001001010101001011001 ;
        92:  q   <=  32'b10111111011001100000111110000111 ;
        93:  q   <=  32'b10111111011001110110101111010111 ;
        94:  q   <=  32'b10111111011010001011111100111011 ;
        95:  q   <=  32'b10111111011010100000100110100110 ;
        96:  q   <=  32'b10111111011010110100101100001011 ;
        97:  q   <=  32'b10111111011011001000001101011110 ;
        98:  q   <=  32'b10111111011011011011001010010011 ;
        99:  q   <=  32'b10111111011011101101100010011101 ;
        100:  q   <=  32'b10111111011011111111010101110011 ;
        101:  q   <=  32'b10111111011100010000100100001000 ;
        102:  q   <=  32'b10111111011100100001001101010010 ;
        103:  q   <=  32'b10111111011100110001010001000111 ;
        104:  q   <=  32'b10111111011101000000101111011101 ;
        105:  q   <=  32'b10111111011101001111101000001010 ;
        106:  q   <=  32'b10111111011101011101111011000110 ;
        107:  q   <=  32'b10111111011101101011101000000111 ;
        108:  q   <=  32'b10111111011101111000101111000101 ;
        109:  q   <=  32'b10111111011110000101001111110111 ;
        110:  q   <=  32'b10111111011110010001001010010111 ;
        111:  q   <=  32'b10111111011110011100011110011101 ;
        112:  q   <=  32'b10111111011110100111001100000001 ;
        113:  q   <=  32'b10111111011110110001010010111110 ;
        114:  q   <=  32'b10111111011110111010110011001101 ;
        115:  q   <=  32'b10111111011111000011101100100111 ;
        116:  q   <=  32'b10111111011111001011111111001001 ;
        117:  q   <=  32'b10111111011111010011101010101011 ;
        118:  q   <=  32'b10111111011111011010101111001011 ;
        119:  q   <=  32'b10111111011111100001001100100011 ;
        120:  q   <=  32'b10111111011111100111000010101111 ;
        121:  q   <=  32'b10111111011111101100010001101101 ;
        122:  q   <=  32'b10111111011111110000111001010111 ;
        123:  q   <=  32'b10111111011111110100111001101101 ;
        124:  q   <=  32'b10111111011111111000010010101011 ;
        125:  q   <=  32'b10111111011111111011000100001111 ;
        126:  q   <=  32'b10111111011111111101001110010111 ;
        127:  q   <=  32'b10111111011111111110110001000011 ;
        128:  q   <=  32'b10111111011111111111101100010000 ;
        129:  q   <=  32'b10111111100000000000000000000000 ;
        130:  q   <=  32'b10111111011111111111101100010000 ;
        131:  q   <=  32'b10111111011111111110110001000011 ;
        132:  q   <=  32'b10111111011111111101001110010111 ;
        133:  q   <=  32'b10111111011111111011000100001111 ;
        134:  q   <=  32'b10111111011111111000010010101011 ;
        135:  q   <=  32'b10111111011111110100111001101101 ;
        136:  q   <=  32'b10111111011111110000111001010111 ;
        137:  q   <=  32'b10111111011111101100010001101101 ;
        138:  q   <=  32'b10111111011111100111000010101111 ;
        139:  q   <=  32'b10111111011111100001001100100011 ;
        140:  q   <=  32'b10111111011111011010101111001011 ;
        141:  q   <=  32'b10111111011111010011101010101011 ;
        142:  q   <=  32'b10111111011111001011111111001001 ;
        143:  q   <=  32'b10111111011111000011101100100111 ;
        144:  q   <=  32'b10111111011110111010110011001101 ;
        145:  q   <=  32'b10111111011110110001010010111110 ;
        146:  q   <=  32'b10111111011110100111001100000001 ;
        147:  q   <=  32'b10111111011110011100011110011101 ;
        148:  q   <=  32'b10111111011110010001001010010111 ;
        149:  q   <=  32'b10111111011110000101001111110111 ;
        150:  q   <=  32'b10111111011101111000101111000101 ;
        151:  q   <=  32'b10111111011101101011101000000111 ;
        152:  q   <=  32'b10111111011101011101111011000110 ;
        153:  q   <=  32'b10111111011101001111101000001010 ;
        154:  q   <=  32'b10111111011101000000101111011101 ;
        155:  q   <=  32'b10111111011100110001010001000111 ;
        156:  q   <=  32'b10111111011100100001001101010010 ;
        157:  q   <=  32'b10111111011100010000100100001000 ;
        158:  q   <=  32'b10111111011011111111010101110011 ;
        159:  q   <=  32'b10111111011011101101100010011101 ;
        160:  q   <=  32'b10111111011011011011001010010011 ;
        161:  q   <=  32'b10111111011011001000001101011110 ;
        162:  q   <=  32'b10111111011010110100101100001011 ;
        163:  q   <=  32'b10111111011010100000100110100110 ;
        164:  q   <=  32'b10111111011010001011111100111011 ;
        165:  q   <=  32'b10111111011001110110101111010111 ;
        166:  q   <=  32'b10111111011001100000111110000111 ;
        167:  q   <=  32'b10111111011001001010101001011001 ;
        168:  q   <=  32'b10111111011000110011110001011001 ;
        169:  q   <=  32'b10111111011000011100010110010111 ;
        170:  q   <=  32'b10111111011000000100011000100001 ;
        171:  q   <=  32'b10111111010111101011111000000101 ;
        172:  q   <=  32'b10111111010111010010110101010011 ;
        173:  q   <=  32'b10111111010110111001010000011010 ;
        174:  q   <=  32'b10111111010110011111001001101001 ;
        175:  q   <=  32'b10111111010110000100100001010010 ;
        176:  q   <=  32'b10111111010101101001010111100100 ;
        177:  q   <=  32'b10111111010101001101101100110001 ;
        178:  q   <=  32'b10111111010100110001100001001000 ;
        179:  q   <=  32'b10111111010100010100110100111101 ;
        180:  q   <=  32'b10111111010011110111101000011111 ;
        181:  q   <=  32'b10111111010011011001111100000010 ;
        182:  q   <=  32'b10111111010010111011101111110111 ;
        183:  q   <=  32'b10111111010010011101000100010010 ;
        184:  q   <=  32'b10111111010001111101111001100101 ;
        185:  q   <=  32'b10111111010001011110010000000011 ;
        186:  q   <=  32'b10111111010000111110001000000000 ;
        187:  q   <=  32'b10111111010000011101100001110000 ;
        188:  q   <=  32'b10111111001111111100011101100111 ;
        189:  q   <=  32'b10111111001111011010111011111001 ;
        190:  q   <=  32'b10111111001110111000111100111010 ;
        191:  q   <=  32'b10111111001110010110100001000001 ;
        192:  q   <=  32'b10111111001101110011101000100010 ;
        193:  q   <=  32'b10111111001101010000010011110011 ;
        194:  q   <=  32'b10111111001100101100100011001001 ;
        195:  q   <=  32'b10111111001100001000010110111010 ;
        196:  q   <=  32'b10111111001011100011101111011101 ;
        197:  q   <=  32'b10111111001010111110101101001001 ;
        198:  q   <=  32'b10111111001010011001010000010100 ;
        199:  q   <=  32'b10111111001001110011011001010101 ;
        200:  q   <=  32'b10111111001001001101001000100100 ;
        201:  q   <=  32'b10111111001000100110011110011001 ;
        202:  q   <=  32'b10111111000111111111011011001010 ;
        203:  q   <=  32'b10111111000111010111111111010001 ;
        204:  q   <=  32'b10111111000110110000001011000101 ;
        205:  q   <=  32'b10111111000110000111111110111111 ;
        206:  q   <=  32'b10111111000101011111011011011001 ;
        207:  q   <=  32'b10111111000100110110100000101010 ;
        208:  q   <=  32'b10111111000100001101001111001100 ;
        209:  q   <=  32'b10111111000011100011100111011001 ;
        210:  q   <=  32'b10111111000010111001101001101011 ;
        211:  q   <=  32'b10111111000010001111010110011010 ;
        212:  q   <=  32'b10111111000001100100101110000010 ;
        213:  q   <=  32'b10111111000000111001110000111100 ;
        214:  q   <=  32'b10111111000000001110011111100100 ;
        215:  q   <=  32'b10111110111111000101110100100110 ;
        216:  q   <=  32'b10111110111101101110000011001010 ;
        217:  q   <=  32'b10111110111100010101101011101001 ;
        218:  q   <=  32'b10111110111010111100101110111010 ;
        219:  q   <=  32'b10111110111001100011001101110100 ;
        220:  q   <=  32'b10111110111000001001001001001110 ;
        221:  q   <=  32'b10111110110110101110100010000000 ;
        222:  q   <=  32'b10111110110101010011011001000001 ;
        223:  q   <=  32'b10111110110011110111101111001010 ;
        224:  q   <=  32'b10111110110010011011100101010011 ;
        225:  q   <=  32'b10111110110000111110111100010101 ;
        226:  q   <=  32'b10111110101111100001110101001001 ;
        227:  q   <=  32'b10111110101110000100010000101001 ;
        228:  q   <=  32'b10111110101100100110001111101110 ;
        229:  q   <=  32'b10111110101011000111110011010011 ;
        230:  q   <=  32'b10111110101001101000111100010010 ;
        231:  q   <=  32'b10111110101000001001101011100100 ;
        232:  q   <=  32'b10111110100110101010000010000110 ;
        233:  q   <=  32'b10111110100101001010000000110001 ;
        234:  q   <=  32'b10111110100011101001101000100001 ;
        235:  q   <=  32'b10111110100010001000111010010011 ;
        236:  q   <=  32'b10111110100000100111110111000000 ;
        237:  q   <=  32'b10111110011110001100111111001011 ;
        238:  q   <=  32'b10111110011011001001101001111111 ;
        239:  q   <=  32'b10111110011000000101110000010011 ;
        240:  q   <=  32'b10111110010101000001010100000001 ;
        241:  q   <=  32'b10111110010001111100010111000001 ;
        242:  q   <=  32'b10111110001110110110111011001110 ;
        243:  q   <=  32'b10111110001011110001000010100010 ;
        244:  q   <=  32'b10111110001000101010101110110101 ;
        245:  q   <=  32'b10111110000101100100000010000011 ;
        246:  q   <=  32'b10111110000010011100111110000110 ;
        247:  q   <=  32'b10111101111110101011001001110010 ;
        248:  q   <=  32'b10111101111000011011110000101110 ;
        249:  q   <=  32'b10111101110010001011110100110101 ;
        250:  q   <=  32'b10111101101011111011011010000000 ;
        251:  q   <=  32'b10111101100101101010100100000100 ;
        252:  q   <=  32'b10111101011110110010101101110011 ;
        253:  q   <=  32'b10111101010010001111101100101111 ;
        254:  q   <=  32'b10111101000101101100001100101011 ;
        255:  q   <=  32'b10111100110010010000101010101111 ;
        256:  q   <=  32'b10111100010010010000111010001111 ;
        257:  q   <=  32'b10100101000011010011000100110001 ;
        258:  q   <=  32'b00111100010010010000111010001111 ;
        259:  q   <=  32'b00111100110010010000101010101111 ;
        260:  q   <=  32'b00111101000101101100001100101011 ;
        261:  q   <=  32'b00111101010010001111101100101111 ;
        262:  q   <=  32'b00111101011110110010101101110011 ;
        263:  q   <=  32'b00111101100101101010100100000100 ;
        264:  q   <=  32'b00111101101011111011011010000000 ;
        265:  q   <=  32'b00111101110010001011110100110101 ;
        266:  q   <=  32'b00111101111000011011110000101110 ;
        267:  q   <=  32'b00111101111110101011001001110010 ;
        268:  q   <=  32'b00111110000010011100111110000110 ;
        269:  q   <=  32'b00111110000101100100000010000011 ;
        270:  q   <=  32'b00111110001000101010101110110101 ;
        271:  q   <=  32'b00111110001011110001000010100010 ;
        272:  q   <=  32'b00111110001110110110111011001110 ;
        273:  q   <=  32'b00111110010001111100010111000001 ;
        274:  q   <=  32'b00111110010101000001010100000001 ;
        275:  q   <=  32'b00111110011000000101110000010011 ;
        276:  q   <=  32'b00111110011011001001101001111111 ;
        277:  q   <=  32'b00111110011110001100111111001011 ;
        278:  q   <=  32'b00111110100000100111110111000000 ;
        279:  q   <=  32'b00111110100010001000111010010011 ;
        280:  q   <=  32'b00111110100011101001101000100001 ;
        281:  q   <=  32'b00111110100101001010000000110001 ;
        282:  q   <=  32'b00111110100110101010000010000110 ;
        283:  q   <=  32'b00111110101000001001101011100100 ;
        284:  q   <=  32'b00111110101001101000111100010010 ;
        285:  q   <=  32'b00111110101011000111110011010011 ;
        286:  q   <=  32'b00111110101100100110001111101110 ;
        287:  q   <=  32'b00111110101110000100010000101001 ;
        288:  q   <=  32'b00111110101111100001110101001001 ;
        289:  q   <=  32'b00111110110000111110111100010101 ;
        290:  q   <=  32'b00111110110010011011100101010011 ;
        291:  q   <=  32'b00111110110011110111101111001010 ;
        292:  q   <=  32'b00111110110101010011011001000001 ;
        293:  q   <=  32'b00111110110110101110100010000000 ;
        294:  q   <=  32'b00111110111000001001001001001110 ;
        295:  q   <=  32'b00111110111001100011001101110100 ;
        296:  q   <=  32'b00111110111010111100101110111010 ;
        297:  q   <=  32'b00111110111100010101101011101001 ;
        298:  q   <=  32'b00111110111101101110000011001010 ;
        299:  q   <=  32'b00111110111111000101110100100110 ;
        300:  q   <=  32'b00111111000000001110011111100100 ;
        301:  q   <=  32'b00111111000000111001110000111100 ;
        302:  q   <=  32'b00111111000001100100101110000010 ;
        303:  q   <=  32'b00111111000010001111010110011010 ;
        304:  q   <=  32'b00111111000010111001101001101011 ;
        305:  q   <=  32'b00111111000011100011100111011001 ;
        306:  q   <=  32'b00111111000100001101001111001100 ;
        307:  q   <=  32'b00111111000100110110100000101010 ;
        308:  q   <=  32'b00111111000101011111011011011001 ;
        309:  q   <=  32'b00111111000110000111111110111111 ;
        310:  q   <=  32'b00111111000110110000001011000101 ;
        311:  q   <=  32'b00111111000111010111111111010001 ;
        312:  q   <=  32'b00111111000111111111011011001010 ;
        313:  q   <=  32'b00111111001000100110011110011001 ;
        314:  q   <=  32'b00111111001001001101001000100100 ;
        315:  q   <=  32'b00111111001001110011011001010101 ;
        316:  q   <=  32'b00111111001010011001010000010100 ;
        317:  q   <=  32'b00111111001010111110101101001001 ;
        318:  q   <=  32'b00111111001011100011101111011101 ;
        319:  q   <=  32'b00111111001100001000010110111010 ;
        320:  q   <=  32'b00111111001100101100100011001001 ;
        321:  q   <=  32'b00111111001101010000010011110011 ;
        322:  q   <=  32'b00111111001101110011101000100010 ;
        323:  q   <=  32'b00111111001110010110100001000001 ;
        324:  q   <=  32'b00111111001110111000111100111010 ;
        325:  q   <=  32'b00111111001111011010111011111001 ;
        326:  q   <=  32'b00111111001111111100011101100111 ;
        327:  q   <=  32'b00111111010000011101100001110000 ;
        328:  q   <=  32'b00111111010000111110001000000000 ;
        329:  q   <=  32'b00111111010001011110010000000011 ;
        330:  q   <=  32'b00111111010001111101111001100101 ;
        331:  q   <=  32'b00111111010010011101000100010010 ;
        332:  q   <=  32'b00111111010010111011101111110111 ;
        333:  q   <=  32'b00111111010011011001111100000010 ;
        334:  q   <=  32'b00111111010011110111101000011111 ;
        335:  q   <=  32'b00111111010100010100110100111101 ;
        336:  q   <=  32'b00111111010100110001100001001000 ;
        337:  q   <=  32'b00111111010101001101101100110001 ;
        338:  q   <=  32'b00111111010101101001010111100100 ;
        339:  q   <=  32'b00111111010110000100100001010010 ;
        340:  q   <=  32'b00111111010110011111001001101001 ;
        341:  q   <=  32'b00111111010110111001010000011010 ;
        342:  q   <=  32'b00111111010111010010110101010011 ;
        343:  q   <=  32'b00111111010111101011111000000101 ;
        344:  q   <=  32'b00111111011000000100011000100001 ;
        345:  q   <=  32'b00111111011000011100010110010111 ;
        346:  q   <=  32'b00111111011000110011110001011001 ;
        347:  q   <=  32'b00111111011001001010101001011001 ;
        348:  q   <=  32'b00111111011001100000111110000111 ;
        349:  q   <=  32'b00111111011001110110101111010111 ;
        350:  q   <=  32'b00111111011010001011111100111011 ;
        351:  q   <=  32'b00111111011010100000100110100110 ;
        352:  q   <=  32'b00111111011010110100101100001011 ;
        353:  q   <=  32'b00111111011011001000001101011110 ;
        354:  q   <=  32'b00111111011011011011001010010011 ;
        355:  q   <=  32'b00111111011011101101100010011101 ;
        356:  q   <=  32'b00111111011011111111010101110011 ;
        357:  q   <=  32'b00111111011100010000100100001000 ;
        358:  q   <=  32'b00111111011100100001001101010010 ;
        359:  q   <=  32'b00111111011100110001010001000111 ;
        360:  q   <=  32'b00111111011101000000101111011101 ;
        361:  q   <=  32'b00111111011101001111101000001010 ;
        362:  q   <=  32'b00111111011101011101111011000110 ;
        363:  q   <=  32'b00111111011101101011101000000111 ;
        364:  q   <=  32'b00111111011101111000101111000101 ;
        365:  q   <=  32'b00111111011110000101001111110111 ;
        366:  q   <=  32'b00111111011110010001001010010111 ;
        367:  q   <=  32'b00111111011110011100011110011101 ;
        368:  q   <=  32'b00111111011110100111001100000001 ;
        369:  q   <=  32'b00111111011110110001010010111110 ;
        370:  q   <=  32'b00111111011110111010110011001101 ;
        371:  q   <=  32'b00111111011111000011101100100111 ;
        372:  q   <=  32'b00111111011111001011111111001001 ;
        373:  q   <=  32'b00111111011111010011101010101011 ;
        374:  q   <=  32'b00111111011111011010101111001011 ;
        375:  q   <=  32'b00111111011111100001001100100011 ;
        376:  q   <=  32'b00111111011111100111000010101111 ;
        377:  q   <=  32'b00111111011111101100010001101101 ;
        378:  q   <=  32'b00111111011111110000111001010111 ;
        379:  q   <=  32'b00111111011111110100111001101101 ;
        380:  q   <=  32'b00111111011111111000010010101011 ;
        381:  q   <=  32'b00111111011111111011000100001111 ;
        382:  q   <=  32'b00111111011111111101001110010111 ;
        383:  q   <=  32'b00111111011111111110110001000011 ;
        384:  q   <=  32'b00111111011111111111101100010000 ;
        385:  q   <=  32'b00111111100000000000000000000000 ;
        386:  q   <=  32'b00111111011111111111101100010000 ;
        387:  q   <=  32'b00111111011111111110110001000011 ;
        388:  q   <=  32'b00111111011111111101001110010111 ;
        389:  q   <=  32'b00111111011111111011000100001111 ;
        390:  q   <=  32'b00111111011111111000010010101011 ;
        391:  q   <=  32'b00111111011111110100111001101101 ;
        392:  q   <=  32'b00111111011111110000111001010111 ;
        393:  q   <=  32'b00111111011111101100010001101101 ;
        394:  q   <=  32'b00111111011111100111000010101111 ;
        395:  q   <=  32'b00111111011111100001001100100011 ;
        396:  q   <=  32'b00111111011111011010101111001011 ;
        397:  q   <=  32'b00111111011111010011101010101011 ;
        398:  q   <=  32'b00111111011111001011111111001001 ;
        399:  q   <=  32'b00111111011111000011101100100111 ;
        400:  q   <=  32'b00111111011110111010110011001101 ;
        401:  q   <=  32'b00111111011110110001010010111110 ;
        402:  q   <=  32'b00111111011110100111001100000001 ;
        403:  q   <=  32'b00111111011110011100011110011101 ;
        404:  q   <=  32'b00111111011110010001001010010111 ;
        405:  q   <=  32'b00111111011110000101001111110111 ;
        406:  q   <=  32'b00111111011101111000101111000101 ;
        407:  q   <=  32'b00111111011101101011101000000111 ;
        408:  q   <=  32'b00111111011101011101111011000110 ;
        409:  q   <=  32'b00111111011101001111101000001010 ;
        410:  q   <=  32'b00111111011101000000101111011101 ;
        411:  q   <=  32'b00111111011100110001010001000111 ;
        412:  q   <=  32'b00111111011100100001001101010010 ;
        413:  q   <=  32'b00111111011100010000100100001000 ;
        414:  q   <=  32'b00111111011011111111010101110011 ;
        415:  q   <=  32'b00111111011011101101100010011101 ;
        416:  q   <=  32'b00111111011011011011001010010011 ;
        417:  q   <=  32'b00111111011011001000001101011110 ;
        418:  q   <=  32'b00111111011010110100101100001011 ;
        419:  q   <=  32'b00111111011010100000100110100110 ;
        420:  q   <=  32'b00111111011010001011111100111011 ;
        421:  q   <=  32'b00111111011001110110101111010111 ;
        422:  q   <=  32'b00111111011001100000111110000111 ;
        423:  q   <=  32'b00111111011001001010101001011001 ;
        424:  q   <=  32'b00111111011000110011110001011001 ;
        425:  q   <=  32'b00111111011000011100010110010111 ;
        426:  q   <=  32'b00111111011000000100011000100001 ;
        427:  q   <=  32'b00111111010111101011111000000101 ;
        428:  q   <=  32'b00111111010111010010110101010011 ;
        429:  q   <=  32'b00111111010110111001010000011010 ;
        430:  q   <=  32'b00111111010110011111001001101001 ;
        431:  q   <=  32'b00111111010110000100100001010010 ;
        432:  q   <=  32'b00111111010101101001010111100100 ;
        433:  q   <=  32'b00111111010101001101101100110001 ;
        434:  q   <=  32'b00111111010100110001100001001000 ;
        435:  q   <=  32'b00111111010100010100110100111101 ;
        436:  q   <=  32'b00111111010011110111101000011111 ;
        437:  q   <=  32'b00111111010011011001111100000010 ;
        438:  q   <=  32'b00111111010010111011101111110111 ;
        439:  q   <=  32'b00111111010010011101000100010010 ;
        440:  q   <=  32'b00111111010001111101111001100101 ;
        441:  q   <=  32'b00111111010001011110010000000011 ;
        442:  q   <=  32'b00111111010000111110001000000000 ;
        443:  q   <=  32'b00111111010000011101100001110000 ;
        444:  q   <=  32'b00111111001111111100011101100111 ;
        445:  q   <=  32'b00111111001111011010111011111001 ;
        446:  q   <=  32'b00111111001110111000111100111010 ;
        447:  q   <=  32'b00111111001110010110100001000001 ;
        448:  q   <=  32'b00111111001101110011101000100010 ;
        449:  q   <=  32'b00111111001101010000010011110011 ;
        450:  q   <=  32'b00111111001100101100100011001001 ;
        451:  q   <=  32'b00111111001100001000010110111010 ;
        452:  q   <=  32'b00111111001011100011101111011101 ;
        453:  q   <=  32'b00111111001010111110101101001001 ;
        454:  q   <=  32'b00111111001010011001010000010100 ;
        455:  q   <=  32'b00111111001001110011011001010101 ;
        456:  q   <=  32'b00111111001001001101001000100100 ;
        457:  q   <=  32'b00111111001000100110011110011001 ;
        458:  q   <=  32'b00111111000111111111011011001010 ;
        459:  q   <=  32'b00111111000111010111111111010001 ;
        460:  q   <=  32'b00111111000110110000001011000101 ;
        461:  q   <=  32'b00111111000110000111111110111111 ;
        462:  q   <=  32'b00111111000101011111011011011001 ;
        463:  q   <=  32'b00111111000100110110100000101010 ;
        464:  q   <=  32'b00111111000100001101001111001100 ;
        465:  q   <=  32'b00111111000011100011100111011001 ;
        466:  q   <=  32'b00111111000010111001101001101011 ;
        467:  q   <=  32'b00111111000010001111010110011010 ;
        468:  q   <=  32'b00111111000001100100101110000010 ;
        469:  q   <=  32'b00111111000000111001110000111100 ;
        470:  q   <=  32'b00111111000000001110011111100100 ;
        471:  q   <=  32'b00111110111111000101110100100110 ;
        472:  q   <=  32'b00111110111101101110000011001010 ;
        473:  q   <=  32'b00111110111100010101101011101001 ;
        474:  q   <=  32'b00111110111010111100101110111010 ;
        475:  q   <=  32'b00111110111001100011001101110100 ;
        476:  q   <=  32'b00111110111000001001001001001110 ;
        477:  q   <=  32'b00111110110110101110100010000000 ;
        478:  q   <=  32'b00111110110101010011011001000001 ;
        479:  q   <=  32'b00111110110011110111101111001010 ;
        480:  q   <=  32'b00111110110010011011100101010011 ;
        481:  q   <=  32'b00111110110000111110111100010101 ;
        482:  q   <=  32'b00111110101111100001110101001001 ;
        483:  q   <=  32'b00111110101110000100010000101001 ;
        484:  q   <=  32'b00111110101100100110001111101110 ;
        485:  q   <=  32'b00111110101011000111110011010011 ;
        486:  q   <=  32'b00111110101001101000111100010010 ;
        487:  q   <=  32'b00111110101000001001101011100100 ;
        488:  q   <=  32'b00111110100110101010000010000110 ;
        489:  q   <=  32'b00111110100101001010000000110001 ;
        490:  q   <=  32'b00111110100011101001101000100001 ;
        491:  q   <=  32'b00111110100010001000111010010011 ;
        492:  q   <=  32'b00111110100000100111110111000000 ;
        493:  q   <=  32'b00111110011110001100111111001011 ;
        494:  q   <=  32'b00111110011011001001101001111111 ;
        495:  q   <=  32'b00111110011000000101110000010011 ;
        496:  q   <=  32'b00111110010101000001010100000001 ;
        497:  q   <=  32'b00111110010001111100010111000001 ;
        498:  q   <=  32'b00111110001110110110111011001110 ;
        499:  q   <=  32'b00111110001011110001000010100010 ;
        500:  q   <=  32'b00111110001000101010101110110101 ;
        501:  q   <=  32'b00111110000101100100000010000011 ;
        502:  q   <=  32'b00111110000010011100111110000110 ;
        503:  q   <=  32'b00111101111110101011001001110010 ;
        504:  q   <=  32'b00111101111000011011110000101110 ;
        505:  q   <=  32'b00111101110010001011110100110101 ;
        506:  q   <=  32'b00111101101011111011011010000000 ;
        507:  q   <=  32'b00111101100101101010100100000100 ;
        508:  q   <=  32'b00111101011110110010101101110011 ;
        509:  q   <=  32'b00111101010010001111101100101111 ;
        510:  q   <=  32'b00111101000101101100001100101011 ;
        511:  q   <=  32'b00111100110010010000101010101111 ;
        512:  q   <=  32'b00111100010010010000111010001111;
        default: q <= 0;
    endcase
end
endmodule
