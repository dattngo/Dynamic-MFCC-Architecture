module mem_w_real (clk, addr, cen, wen, data,q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00111111100000000000000000000000 ;
        2:  q   <=  32'b00111111011111111111101100010000 ;
        3:  q   <=  32'b00111111011111111110110001000011 ;
        4:  q   <=  32'b00111111011111111101001110010111 ;
        5:  q   <=  32'b00111111011111111011000100001111 ;
        6:  q   <=  32'b00111111011111111000010010101011 ;
        7:  q   <=  32'b00111111011111110100111001101101 ;
        8:  q   <=  32'b00111111011111110000111001010111 ;
        9:  q   <=  32'b00111111011111101100010001101101 ;
        10:  q   <=  32'b00111111011111100111000010101111 ;
        11:  q   <=  32'b00111111011111100001001100100011 ;
        12:  q   <=  32'b00111111011111011010101111001011 ;
        13:  q   <=  32'b00111111011111010011101010101011 ;
        14:  q   <=  32'b00111111011111001011111111001001 ;
        15:  q   <=  32'b00111111011111000011101100100111 ;
        16:  q   <=  32'b00111111011110111010110011001101 ;
        17:  q   <=  32'b00111111011110110001010010111110 ;
        18:  q   <=  32'b00111111011110100111001100000001 ;
        19:  q   <=  32'b00111111011110011100011110011101 ;
        20:  q   <=  32'b00111111011110010001001010010111 ;
        21:  q   <=  32'b00111111011110000101001111110111 ;
        22:  q   <=  32'b00111111011101111000101111000101 ;
        23:  q   <=  32'b00111111011101101011101000000111 ;
        24:  q   <=  32'b00111111011101011101111011000110 ;
        25:  q   <=  32'b00111111011101001111101000001010 ;
        26:  q   <=  32'b00111111011101000000101111011101 ;
        27:  q   <=  32'b00111111011100110001010001000111 ;
        28:  q   <=  32'b00111111011100100001001101010010 ;
        29:  q   <=  32'b00111111011100010000100100001000 ;
        30:  q   <=  32'b00111111011011111111010101110011 ;
        31:  q   <=  32'b00111111011011101101100010011101 ;
        32:  q   <=  32'b00111111011011011011001010010011 ;
        33:  q   <=  32'b00111111011011001000001101011110 ;
        34:  q   <=  32'b00111111011010110100101100001011 ;
        35:  q   <=  32'b00111111011010100000100110100110 ;
        36:  q   <=  32'b00111111011010001011111100111011 ;
        37:  q   <=  32'b00111111011001110110101111010111 ;
        38:  q   <=  32'b00111111011001100000111110000111 ;
        39:  q   <=  32'b00111111011001001010101001011001 ;
        40:  q   <=  32'b00111111011000110011110001011001 ;
        41:  q   <=  32'b00111111011000011100010110010111 ;
        42:  q   <=  32'b00111111011000000100011000100001 ;
        43:  q   <=  32'b00111111010111101011111000000101 ;
        44:  q   <=  32'b00111111010111010010110101010011 ;
        45:  q   <=  32'b00111111010110111001010000011010 ;
        46:  q   <=  32'b00111111010110011111001001101001 ;
        47:  q   <=  32'b00111111010110000100100001010010 ;
        48:  q   <=  32'b00111111010101101001010111100100 ;
        49:  q   <=  32'b00111111010101001101101100110001 ;
        50:  q   <=  32'b00111111010100110001100001001000 ;
        51:  q   <=  32'b00111111010100010100110100111101 ;
        52:  q   <=  32'b00111111010011110111101000011111 ;
        53:  q   <=  32'b00111111010011011001111100000010 ;
        54:  q   <=  32'b00111111010010111011101111110111 ;
        55:  q   <=  32'b00111111010010011101000100010010 ;
        56:  q   <=  32'b00111111010001111101111001100101 ;
        57:  q   <=  32'b00111111010001011110010000000011 ;
        58:  q   <=  32'b00111111010000111110001000000000 ;
        59:  q   <=  32'b00111111010000011101100001110000 ;
        60:  q   <=  32'b00111111001111111100011101100111 ;
        61:  q   <=  32'b00111111001111011010111011111001 ;
        62:  q   <=  32'b00111111001110111000111100111010 ;
        63:  q   <=  32'b00111111001110010110100001000001 ;
        64:  q   <=  32'b00111111001101110011101000100010 ;
        65:  q   <=  32'b00111111001101010000010011110011 ;
        66:  q   <=  32'b00111111001100101100100011001001 ;
        67:  q   <=  32'b00111111001100001000010110111010 ;
        68:  q   <=  32'b00111111001011100011101111011101 ;
        69:  q   <=  32'b00111111001010111110101101001001 ;
        70:  q   <=  32'b00111111001010011001010000010100 ;
        71:  q   <=  32'b00111111001001110011011001010101 ;
        72:  q   <=  32'b00111111001001001101001000100100 ;
        73:  q   <=  32'b00111111001000100110011110011001 ;
        74:  q   <=  32'b00111111000111111111011011001010 ;
        75:  q   <=  32'b00111111000111010111111111010001 ;
        76:  q   <=  32'b00111111000110110000001011000101 ;
        77:  q   <=  32'b00111111000110000111111110111111 ;
        78:  q   <=  32'b00111111000101011111011011011001 ;
        79:  q   <=  32'b00111111000100110110100000101010 ;
        80:  q   <=  32'b00111111000100001101001111001100 ;
        81:  q   <=  32'b00111111000011100011100111011001 ;
        82:  q   <=  32'b00111111000010111001101001101011 ;
        83:  q   <=  32'b00111111000010001111010110011010 ;
        84:  q   <=  32'b00111111000001100100101110000010 ;
        85:  q   <=  32'b00111111000000111001110000111100 ;
        86:  q   <=  32'b00111111000000001110011111100100 ;
        87:  q   <=  32'b00111110111111000101110100100110 ;
        88:  q   <=  32'b00111110111101101110000011001010 ;
        89:  q   <=  32'b00111110111100010101101011101001 ;
        90:  q   <=  32'b00111110111010111100101110111010 ;
        91:  q   <=  32'b00111110111001100011001101110100 ;
        92:  q   <=  32'b00111110111000001001001001001110 ;
        93:  q   <=  32'b00111110110110101110100010000000 ;
        94:  q   <=  32'b00111110110101010011011001000001 ;
        95:  q   <=  32'b00111110110011110111101111001010 ;
        96:  q   <=  32'b00111110110010011011100101010011 ;
        97:  q   <=  32'b00111110110000111110111100010101 ;
        98:  q   <=  32'b00111110101111100001110101001001 ;
        99:  q   <=  32'b00111110101110000100010000101001 ;
        100:  q   <=  32'b00111110101100100110001111101110 ;
        101:  q   <=  32'b00111110101011000111110011010011 ;
        102:  q   <=  32'b00111110101001101000111100010010 ;
        103:  q   <=  32'b00111110101000001001101011100100 ;
        104:  q   <=  32'b00111110100110101010000010000110 ;
        105:  q   <=  32'b00111110100101001010000000110001 ;
        106:  q   <=  32'b00111110100011101001101000100001 ;
        107:  q   <=  32'b00111110100010001000111010010011 ;
        108:  q   <=  32'b00111110100000100111110111000000 ;
        109:  q   <=  32'b00111110011110001100111111001011 ;
        110:  q   <=  32'b00111110011011001001101001111111 ;
        111:  q   <=  32'b00111110011000000101110000010011 ;
        112:  q   <=  32'b00111110010101000001010100000001 ;
        113:  q   <=  32'b00111110010001111100010111000001 ;
        114:  q   <=  32'b00111110001110110110111011001110 ;
        115:  q   <=  32'b00111110001011110001000010100010 ;
        116:  q   <=  32'b00111110001000101010101110110101 ;
        117:  q   <=  32'b00111110000101100100000010000011 ;
        118:  q   <=  32'b00111110000010011100111110000110 ;
        119:  q   <=  32'b00111101111110101011001001110010 ;
        120:  q   <=  32'b00111101111000011011110000101110 ;
        121:  q   <=  32'b00111101110010001011110100110101 ;
        122:  q   <=  32'b00111101101011111011011010000000 ;
        123:  q   <=  32'b00111101100101101010100100000100 ;
        124:  q   <=  32'b00111101011110110010101101110011 ;
        125:  q   <=  32'b00111101010010001111101100101111 ;
        126:  q   <=  32'b00111101000101101100001100101011 ;
        127:  q   <=  32'b00111100110010010000101010101111 ;
        128:  q   <=  32'b00111100010010010000111010001111 ;
        129:  q   <=  32'b00100100100011010011000100110001 ;
        130:  q   <=  32'b10111100010010010000111010001111 ;
        131:  q   <=  32'b10111100110010010000101010101111 ;
        132:  q   <=  32'b10111101000101101100001100101011 ;
        133:  q   <=  32'b10111101010010001111101100101111 ;
        134:  q   <=  32'b10111101011110110010101101110011 ;
        135:  q   <=  32'b10111101100101101010100100000100 ;
        136:  q   <=  32'b10111101101011111011011010000000 ;
        137:  q   <=  32'b10111101110010001011110100110101 ;
        138:  q   <=  32'b10111101111000011011110000101110 ;
        139:  q   <=  32'b10111101111110101011001001110010 ;
        140:  q   <=  32'b10111110000010011100111110000110 ;
        141:  q   <=  32'b10111110000101100100000010000011 ;
        142:  q   <=  32'b10111110001000101010101110110101 ;
        143:  q   <=  32'b10111110001011110001000010100010 ;
        144:  q   <=  32'b10111110001110110110111011001110 ;
        145:  q   <=  32'b10111110010001111100010111000001 ;
        146:  q   <=  32'b10111110010101000001010100000001 ;
        147:  q   <=  32'b10111110011000000101110000010011 ;
        148:  q   <=  32'b10111110011011001001101001111111 ;
        149:  q   <=  32'b10111110011110001100111111001011 ;
        150:  q   <=  32'b10111110100000100111110111000000 ;
        151:  q   <=  32'b10111110100010001000111010010011 ;
        152:  q   <=  32'b10111110100011101001101000100001 ;
        153:  q   <=  32'b10111110100101001010000000110001 ;
        154:  q   <=  32'b10111110100110101010000010000110 ;
        155:  q   <=  32'b10111110101000001001101011100100 ;
        156:  q   <=  32'b10111110101001101000111100010010 ;
        157:  q   <=  32'b10111110101011000111110011010011 ;
        158:  q   <=  32'b10111110101100100110001111101110 ;
        159:  q   <=  32'b10111110101110000100010000101001 ;
        160:  q   <=  32'b10111110101111100001110101001001 ;
        161:  q   <=  32'b10111110110000111110111100010101 ;
        162:  q   <=  32'b10111110110010011011100101010011 ;
        163:  q   <=  32'b10111110110011110111101111001010 ;
        164:  q   <=  32'b10111110110101010011011001000001 ;
        165:  q   <=  32'b10111110110110101110100010000000 ;
        166:  q   <=  32'b10111110111000001001001001001110 ;
        167:  q   <=  32'b10111110111001100011001101110100 ;
        168:  q   <=  32'b10111110111010111100101110111010 ;
        169:  q   <=  32'b10111110111100010101101011101001 ;
        170:  q   <=  32'b10111110111101101110000011001010 ;
        171:  q   <=  32'b10111110111111000101110100100110 ;
        172:  q   <=  32'b10111111000000001110011111100100 ;
        173:  q   <=  32'b10111111000000111001110000111100 ;
        174:  q   <=  32'b10111111000001100100101110000010 ;
        175:  q   <=  32'b10111111000010001111010110011010 ;
        176:  q   <=  32'b10111111000010111001101001101011 ;
        177:  q   <=  32'b10111111000011100011100111011001 ;
        178:  q   <=  32'b10111111000100001101001111001100 ;
        179:  q   <=  32'b10111111000100110110100000101010 ;
        180:  q   <=  32'b10111111000101011111011011011001 ;
        181:  q   <=  32'b10111111000110000111111110111111 ;
        182:  q   <=  32'b10111111000110110000001011000101 ;
        183:  q   <=  32'b10111111000111010111111111010001 ;
        184:  q   <=  32'b10111111000111111111011011001010 ;
        185:  q   <=  32'b10111111001000100110011110011001 ;
        186:  q   <=  32'b10111111001001001101001000100100 ;
        187:  q   <=  32'b10111111001001110011011001010101 ;
        188:  q   <=  32'b10111111001010011001010000010100 ;
        189:  q   <=  32'b10111111001010111110101101001001 ;
        190:  q   <=  32'b10111111001011100011101111011101 ;
        191:  q   <=  32'b10111111001100001000010110111010 ;
        192:  q   <=  32'b10111111001100101100100011001001 ;
        193:  q   <=  32'b10111111001101010000010011110011 ;
        194:  q   <=  32'b10111111001101110011101000100010 ;
        195:  q   <=  32'b10111111001110010110100001000001 ;
        196:  q   <=  32'b10111111001110111000111100111010 ;
        197:  q   <=  32'b10111111001111011010111011111001 ;
        198:  q   <=  32'b10111111001111111100011101100111 ;
        199:  q   <=  32'b10111111010000011101100001110000 ;
        200:  q   <=  32'b10111111010000111110001000000000 ;
        201:  q   <=  32'b10111111010001011110010000000011 ;
        202:  q   <=  32'b10111111010001111101111001100101 ;
        203:  q   <=  32'b10111111010010011101000100010010 ;
        204:  q   <=  32'b10111111010010111011101111110111 ;
        205:  q   <=  32'b10111111010011011001111100000010 ;
        206:  q   <=  32'b10111111010011110111101000011111 ;
        207:  q   <=  32'b10111111010100010100110100111101 ;
        208:  q   <=  32'b10111111010100110001100001001000 ;
        209:  q   <=  32'b10111111010101001101101100110001 ;
        210:  q   <=  32'b10111111010101101001010111100100 ;
        211:  q   <=  32'b10111111010110000100100001010010 ;
        212:  q   <=  32'b10111111010110011111001001101001 ;
        213:  q   <=  32'b10111111010110111001010000011010 ;
        214:  q   <=  32'b10111111010111010010110101010011 ;
        215:  q   <=  32'b10111111010111101011111000000101 ;
        216:  q   <=  32'b10111111011000000100011000100001 ;
        217:  q   <=  32'b10111111011000011100010110010111 ;
        218:  q   <=  32'b10111111011000110011110001011001 ;
        219:  q   <=  32'b10111111011001001010101001011001 ;
        220:  q   <=  32'b10111111011001100000111110000111 ;
        221:  q   <=  32'b10111111011001110110101111010111 ;
        222:  q   <=  32'b10111111011010001011111100111011 ;
        223:  q   <=  32'b10111111011010100000100110100110 ;
        224:  q   <=  32'b10111111011010110100101100001011 ;
        225:  q   <=  32'b10111111011011001000001101011110 ;
        226:  q   <=  32'b10111111011011011011001010010011 ;
        227:  q   <=  32'b10111111011011101101100010011101 ;
        228:  q   <=  32'b10111111011011111111010101110011 ;
        229:  q   <=  32'b10111111011100010000100100001000 ;
        230:  q   <=  32'b10111111011100100001001101010010 ;
        231:  q   <=  32'b10111111011100110001010001000111 ;
        232:  q   <=  32'b10111111011101000000101111011101 ;
        233:  q   <=  32'b10111111011101001111101000001010 ;
        234:  q   <=  32'b10111111011101011101111011000110 ;
        235:  q   <=  32'b10111111011101101011101000000111 ;
        236:  q   <=  32'b10111111011101111000101111000101 ;
        237:  q   <=  32'b10111111011110000101001111110111 ;
        238:  q   <=  32'b10111111011110010001001010010111 ;
        239:  q   <=  32'b10111111011110011100011110011101 ;
        240:  q   <=  32'b10111111011110100111001100000001 ;
        241:  q   <=  32'b10111111011110110001010010111110 ;
        242:  q   <=  32'b10111111011110111010110011001101 ;
        243:  q   <=  32'b10111111011111000011101100100111 ;
        244:  q   <=  32'b10111111011111001011111111001001 ;
        245:  q   <=  32'b10111111011111010011101010101011 ;
        246:  q   <=  32'b10111111011111011010101111001011 ;
        247:  q   <=  32'b10111111011111100001001100100011 ;
        248:  q   <=  32'b10111111011111100111000010101111 ;
        249:  q   <=  32'b10111111011111101100010001101101 ;
        250:  q   <=  32'b10111111011111110000111001010111 ;
        251:  q   <=  32'b10111111011111110100111001101101 ;
        252:  q   <=  32'b10111111011111111000010010101011 ;
        253:  q   <=  32'b10111111011111111011000100001111 ;
        254:  q   <=  32'b10111111011111111101001110010111 ;
        255:  q   <=  32'b10111111011111111110110001000011 ;
        256:  q   <=  32'b10111111011111111111101100010000 ;
        257:  q   <=  32'b10111111100000000000000000000000 ;
        258:  q   <=  32'b10111111011111111111101100010000 ;
        259:  q   <=  32'b10111111011111111110110001000011 ;
        260:  q   <=  32'b10111111011111111101001110010111 ;
        261:  q   <=  32'b10111111011111111011000100001111 ;
        262:  q   <=  32'b10111111011111111000010010101011 ;
        263:  q   <=  32'b10111111011111110100111001101101 ;
        264:  q   <=  32'b10111111011111110000111001010111 ;
        265:  q   <=  32'b10111111011111101100010001101101 ;
        266:  q   <=  32'b10111111011111100111000010101111 ;
        267:  q   <=  32'b10111111011111100001001100100011 ;
        268:  q   <=  32'b10111111011111011010101111001011 ;
        269:  q   <=  32'b10111111011111010011101010101011 ;
        270:  q   <=  32'b10111111011111001011111111001001 ;
        271:  q   <=  32'b10111111011111000011101100100111 ;
        272:  q   <=  32'b10111111011110111010110011001101 ;
        273:  q   <=  32'b10111111011110110001010010111110 ;
        274:  q   <=  32'b10111111011110100111001100000001 ;
        275:  q   <=  32'b10111111011110011100011110011101 ;
        276:  q   <=  32'b10111111011110010001001010010111 ;
        277:  q   <=  32'b10111111011110000101001111110111 ;
        278:  q   <=  32'b10111111011101111000101111000101 ;
        279:  q   <=  32'b10111111011101101011101000000111 ;
        280:  q   <=  32'b10111111011101011101111011000110 ;
        281:  q   <=  32'b10111111011101001111101000001010 ;
        282:  q   <=  32'b10111111011101000000101111011101 ;
        283:  q   <=  32'b10111111011100110001010001000111 ;
        284:  q   <=  32'b10111111011100100001001101010010 ;
        285:  q   <=  32'b10111111011100010000100100001000 ;
        286:  q   <=  32'b10111111011011111111010101110011 ;
        287:  q   <=  32'b10111111011011101101100010011101 ;
        288:  q   <=  32'b10111111011011011011001010010011 ;
        289:  q   <=  32'b10111111011011001000001101011110 ;
        290:  q   <=  32'b10111111011010110100101100001011 ;
        291:  q   <=  32'b10111111011010100000100110100110 ;
        292:  q   <=  32'b10111111011010001011111100111011 ;
        293:  q   <=  32'b10111111011001110110101111010111 ;
        294:  q   <=  32'b10111111011001100000111110000111 ;
        295:  q   <=  32'b10111111011001001010101001011001 ;
        296:  q   <=  32'b10111111011000110011110001011001 ;
        297:  q   <=  32'b10111111011000011100010110010111 ;
        298:  q   <=  32'b10111111011000000100011000100001 ;
        299:  q   <=  32'b10111111010111101011111000000101 ;
        300:  q   <=  32'b10111111010111010010110101010011 ;
        301:  q   <=  32'b10111111010110111001010000011010 ;
        302:  q   <=  32'b10111111010110011111001001101001 ;
        303:  q   <=  32'b10111111010110000100100001010010 ;
        304:  q   <=  32'b10111111010101101001010111100100 ;
        305:  q   <=  32'b10111111010101001101101100110001 ;
        306:  q   <=  32'b10111111010100110001100001001000 ;
        307:  q   <=  32'b10111111010100010100110100111101 ;
        308:  q   <=  32'b10111111010011110111101000011111 ;
        309:  q   <=  32'b10111111010011011001111100000010 ;
        310:  q   <=  32'b10111111010010111011101111110111 ;
        311:  q   <=  32'b10111111010010011101000100010010 ;
        312:  q   <=  32'b10111111010001111101111001100101 ;
        313:  q   <=  32'b10111111010001011110010000000011 ;
        314:  q   <=  32'b10111111010000111110001000000000 ;
        315:  q   <=  32'b10111111010000011101100001110000 ;
        316:  q   <=  32'b10111111001111111100011101100111 ;
        317:  q   <=  32'b10111111001111011010111011111001 ;
        318:  q   <=  32'b10111111001110111000111100111010 ;
        319:  q   <=  32'b10111111001110010110100001000001 ;
        320:  q   <=  32'b10111111001101110011101000100010 ;
        321:  q   <=  32'b10111111001101010000010011110011 ;
        322:  q   <=  32'b10111111001100101100100011001001 ;
        323:  q   <=  32'b10111111001100001000010110111010 ;
        324:  q   <=  32'b10111111001011100011101111011101 ;
        325:  q   <=  32'b10111111001010111110101101001001 ;
        326:  q   <=  32'b10111111001010011001010000010100 ;
        327:  q   <=  32'b10111111001001110011011001010101 ;
        328:  q   <=  32'b10111111001001001101001000100100 ;
        329:  q   <=  32'b10111111001000100110011110011001 ;
        330:  q   <=  32'b10111111000111111111011011001010 ;
        331:  q   <=  32'b10111111000111010111111111010001 ;
        332:  q   <=  32'b10111111000110110000001011000101 ;
        333:  q   <=  32'b10111111000110000111111110111111 ;
        334:  q   <=  32'b10111111000101011111011011011001 ;
        335:  q   <=  32'b10111111000100110110100000101010 ;
        336:  q   <=  32'b10111111000100001101001111001100 ;
        337:  q   <=  32'b10111111000011100011100111011001 ;
        338:  q   <=  32'b10111111000010111001101001101011 ;
        339:  q   <=  32'b10111111000010001111010110011010 ;
        340:  q   <=  32'b10111111000001100100101110000010 ;
        341:  q   <=  32'b10111111000000111001110000111100 ;
        342:  q   <=  32'b10111111000000001110011111100100 ;
        343:  q   <=  32'b10111110111111000101110100100110 ;
        344:  q   <=  32'b10111110111101101110000011001010 ;
        345:  q   <=  32'b10111110111100010101101011101001 ;
        346:  q   <=  32'b10111110111010111100101110111010 ;
        347:  q   <=  32'b10111110111001100011001101110100 ;
        348:  q   <=  32'b10111110111000001001001001001110 ;
        349:  q   <=  32'b10111110110110101110100010000000 ;
        350:  q   <=  32'b10111110110101010011011001000001 ;
        351:  q   <=  32'b10111110110011110111101111001010 ;
        352:  q   <=  32'b10111110110010011011100101010011 ;
        353:  q   <=  32'b10111110110000111110111100010101 ;
        354:  q   <=  32'b10111110101111100001110101001001 ;
        355:  q   <=  32'b10111110101110000100010000101001 ;
        356:  q   <=  32'b10111110101100100110001111101110 ;
        357:  q   <=  32'b10111110101011000111110011010011 ;
        358:  q   <=  32'b10111110101001101000111100010010 ;
        359:  q   <=  32'b10111110101000001001101011100100 ;
        360:  q   <=  32'b10111110100110101010000010000110 ;
        361:  q   <=  32'b10111110100101001010000000110001 ;
        362:  q   <=  32'b10111110100011101001101000100001 ;
        363:  q   <=  32'b10111110100010001000111010010011 ;
        364:  q   <=  32'b10111110100000100111110111000000 ;
        365:  q   <=  32'b10111110011110001100111111001011 ;
        366:  q   <=  32'b10111110011011001001101001111111 ;
        367:  q   <=  32'b10111110011000000101110000010011 ;
        368:  q   <=  32'b10111110010101000001010100000001 ;
        369:  q   <=  32'b10111110010001111100010111000001 ;
        370:  q   <=  32'b10111110001110110110111011001110 ;
        371:  q   <=  32'b10111110001011110001000010100010 ;
        372:  q   <=  32'b10111110001000101010101110110101 ;
        373:  q   <=  32'b10111110000101100100000010000011 ;
        374:  q   <=  32'b10111110000010011100111110000110 ;
        375:  q   <=  32'b10111101111110101011001001110010 ;
        376:  q   <=  32'b10111101111000011011110000101110 ;
        377:  q   <=  32'b10111101110010001011110100110101 ;
        378:  q   <=  32'b10111101101011111011011010000000 ;
        379:  q   <=  32'b10111101100101101010100100000100 ;
        380:  q   <=  32'b10111101011110110010101101110011 ;
        381:  q   <=  32'b10111101010010001111101100101111 ;
        382:  q   <=  32'b10111101000101101100001100101011 ;
        383:  q   <=  32'b10111100110010010000101010101111 ;
        384:  q   <=  32'b10111100010010010000111010001111 ;
        385:  q   <=  32'b10100101010100111100100111001010 ;
        386:  q   <=  32'b00111100010010010000111010001111 ;
        387:  q   <=  32'b00111100110010010000101010101111 ;
        388:  q   <=  32'b00111101000101101100001100101011 ;
        389:  q   <=  32'b00111101010010001111101100101111 ;
        390:  q   <=  32'b00111101011110110010101101110011 ;
        391:  q   <=  32'b00111101100101101010100100000100 ;
        392:  q   <=  32'b00111101101011111011011010000000 ;
        393:  q   <=  32'b00111101110010001011110100110101 ;
        394:  q   <=  32'b00111101111000011011110000101110 ;
        395:  q   <=  32'b00111101111110101011001001110010 ;
        396:  q   <=  32'b00111110000010011100111110000110 ;
        397:  q   <=  32'b00111110000101100100000010000011 ;
        398:  q   <=  32'b00111110001000101010101110110101 ;
        399:  q   <=  32'b00111110001011110001000010100010 ;
        400:  q   <=  32'b00111110001110110110111011001110 ;
        401:  q   <=  32'b00111110010001111100010111000001 ;
        402:  q   <=  32'b00111110010101000001010100000001 ;
        403:  q   <=  32'b00111110011000000101110000010011 ;
        404:  q   <=  32'b00111110011011001001101001111111 ;
        405:  q   <=  32'b00111110011110001100111111001011 ;
        406:  q   <=  32'b00111110100000100111110111000000 ;
        407:  q   <=  32'b00111110100010001000111010010011 ;
        408:  q   <=  32'b00111110100011101001101000100001 ;
        409:  q   <=  32'b00111110100101001010000000110001 ;
        410:  q   <=  32'b00111110100110101010000010000110 ;
        411:  q   <=  32'b00111110101000001001101011100100 ;
        412:  q   <=  32'b00111110101001101000111100010010 ;
        413:  q   <=  32'b00111110101011000111110011010011 ;
        414:  q   <=  32'b00111110101100100110001111101110 ;
        415:  q   <=  32'b00111110101110000100010000101001 ;
        416:  q   <=  32'b00111110101111100001110101001001 ;
        417:  q   <=  32'b00111110110000111110111100010101 ;
        418:  q   <=  32'b00111110110010011011100101010011 ;
        419:  q   <=  32'b00111110110011110111101111001010 ;
        420:  q   <=  32'b00111110110101010011011001000001 ;
        421:  q   <=  32'b00111110110110101110100010000000 ;
        422:  q   <=  32'b00111110111000001001001001001110 ;
        423:  q   <=  32'b00111110111001100011001101110100 ;
        424:  q   <=  32'b00111110111010111100101110111010 ;
        425:  q   <=  32'b00111110111100010101101011101001 ;
        426:  q   <=  32'b00111110111101101110000011001010 ;
        427:  q   <=  32'b00111110111111000101110100100110 ;
        428:  q   <=  32'b00111111000000001110011111100100 ;
        429:  q   <=  32'b00111111000000111001110000111100 ;
        430:  q   <=  32'b00111111000001100100101110000010 ;
        431:  q   <=  32'b00111111000010001111010110011010 ;
        432:  q   <=  32'b00111111000010111001101001101011 ;
        433:  q   <=  32'b00111111000011100011100111011001 ;
        434:  q   <=  32'b00111111000100001101001111001100 ;
        435:  q   <=  32'b00111111000100110110100000101010 ;
        436:  q   <=  32'b00111111000101011111011011011001 ;
        437:  q   <=  32'b00111111000110000111111110111111 ;
        438:  q   <=  32'b00111111000110110000001011000101 ;
        439:  q   <=  32'b00111111000111010111111111010001 ;
        440:  q   <=  32'b00111111000111111111011011001010 ;
        441:  q   <=  32'b00111111001000100110011110011001 ;
        442:  q   <=  32'b00111111001001001101001000100100 ;
        443:  q   <=  32'b00111111001001110011011001010101 ;
        444:  q   <=  32'b00111111001010011001010000010100 ;
        445:  q   <=  32'b00111111001010111110101101001001 ;
        446:  q   <=  32'b00111111001011100011101111011101 ;
        447:  q   <=  32'b00111111001100001000010110111010 ;
        448:  q   <=  32'b00111111001100101100100011001001 ;
        449:  q   <=  32'b00111111001101010000010011110011 ;
        450:  q   <=  32'b00111111001101110011101000100010 ;
        451:  q   <=  32'b00111111001110010110100001000001 ;
        452:  q   <=  32'b00111111001110111000111100111010 ;
        453:  q   <=  32'b00111111001111011010111011111001 ;
        454:  q   <=  32'b00111111001111111100011101100111 ;
        455:  q   <=  32'b00111111010000011101100001110000 ;
        456:  q   <=  32'b00111111010000111110001000000000 ;
        457:  q   <=  32'b00111111010001011110010000000011 ;
        458:  q   <=  32'b00111111010001111101111001100101 ;
        459:  q   <=  32'b00111111010010011101000100010010 ;
        460:  q   <=  32'b00111111010010111011101111110111 ;
        461:  q   <=  32'b00111111010011011001111100000010 ;
        462:  q   <=  32'b00111111010011110111101000011111 ;
        463:  q   <=  32'b00111111010100010100110100111101 ;
        464:  q   <=  32'b00111111010100110001100001001000 ;
        465:  q   <=  32'b00111111010101001101101100110001 ;
        466:  q   <=  32'b00111111010101101001010111100100 ;
        467:  q   <=  32'b00111111010110000100100001010010 ;
        468:  q   <=  32'b00111111010110011111001001101001 ;
        469:  q   <=  32'b00111111010110111001010000011010 ;
        470:  q   <=  32'b00111111010111010010110101010011 ;
        471:  q   <=  32'b00111111010111101011111000000101 ;
        472:  q   <=  32'b00111111011000000100011000100001 ;
        473:  q   <=  32'b00111111011000011100010110010111 ;
        474:  q   <=  32'b00111111011000110011110001011001 ;
        475:  q   <=  32'b00111111011001001010101001011001 ;
        476:  q   <=  32'b00111111011001100000111110000111 ;
        477:  q   <=  32'b00111111011001110110101111010111 ;
        478:  q   <=  32'b00111111011010001011111100111011 ;
        479:  q   <=  32'b00111111011010100000100110100110 ;
        480:  q   <=  32'b00111111011010110100101100001011 ;
        481:  q   <=  32'b00111111011011001000001101011110 ;
        482:  q   <=  32'b00111111011011011011001010010011 ;
        483:  q   <=  32'b00111111011011101101100010011101 ;
        484:  q   <=  32'b00111111011011111111010101110011 ;
        485:  q   <=  32'b00111111011100010000100100001000 ;
        486:  q   <=  32'b00111111011100100001001101010010 ;
        487:  q   <=  32'b00111111011100110001010001000111 ;
        488:  q   <=  32'b00111111011101000000101111011101 ;
        489:  q   <=  32'b00111111011101001111101000001010 ;
        490:  q   <=  32'b00111111011101011101111011000110 ;
        491:  q   <=  32'b00111111011101101011101000000111 ;
        492:  q   <=  32'b00111111011101111000101111000101 ;
        493:  q   <=  32'b00111111011110000101001111110111 ;
        494:  q   <=  32'b00111111011110010001001010010111 ;
        495:  q   <=  32'b00111111011110011100011110011101 ;
        496:  q   <=  32'b00111111011110100111001100000001 ;
        497:  q   <=  32'b00111111011110110001010010111110 ;
        498:  q   <=  32'b00111111011110111010110011001101 ;
        499:  q   <=  32'b00111111011111000011101100100111 ;
        500:  q   <=  32'b00111111011111001011111111001001 ;
        501:  q   <=  32'b00111111011111010011101010101011 ;
        502:  q   <=  32'b00111111011111011010101111001011 ;
        503:  q   <=  32'b00111111011111100001001100100011 ;
        504:  q   <=  32'b00111111011111100111000010101111 ;
        505:  q   <=  32'b00111111011111101100010001101101 ;
        506:  q   <=  32'b00111111011111110000111001010111 ;
        507:  q   <=  32'b00111111011111110100111001101101 ;
        508:  q   <=  32'b00111111011111111000010010101011 ;
        509:  q   <=  32'b00111111011111111011000100001111 ;
        510:  q   <=  32'b00111111011111111101001110010111 ;
        511:  q   <=  32'b00111111011111111110110001000011 ;
        512:  q   <=  32'b00111111011111111111101100010000;
        default: q <= 0;
    endcase
end
endmodule
