module mem_cepstral_cof (clk, addr, cen, wen, data,q);
parameter DATA_WIDTH =  32;
input clk;
input [11:0] addr;
input cen;
input wen;
input [DATA_WIDTH-1:0]data;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clk) begin
    case(addr)
        1:  q   <=  32'b00111111011111111110101110100001 ;
        2:  q   <=  32'b00111111011111110100100010111111 ;
        3:  q   <=  32'b00111111011111100000001101100011 ;
        4:  q   <=  32'b00111111011111000001110001011100 ;
        5:  q   <=  32'b00111111011110011001010011100000 ;
        6:  q   <=  32'b00111111011101100110111010001010 ;
        7:  q   <=  32'b00111111011100101010101101011101 ;
        8:  q   <=  32'b00111111011011100100110110111101 ;
        9:  q   <=  32'b00111111011010010101100001110010 ;
        10:  q   <=  32'b00111111011000111100111010100011 ;
        11:  q   <=  32'b00111111010111011011001111010111 ;
        12:  q   <=  32'b00111111010101110000101111110000 ;
        13:  q   <=  32'b00111111010011111101101100101011 ;
        14:  q   <=  32'b00111111010010000010011000011011 ;
        15:  q   <=  32'b00111111001111111111000110101001 ;
        16:  q   <=  32'b00111111001101110100001100001100 ;
        17:  q   <=  32'b00111111001011100001111111001100 ;
        18:  q   <=  32'b00111111001001001000110110111010 ;
        19:  q   <=  32'b00111111000110101001001011101101 ;
        20:  q   <=  32'b00111111000100000011010110111110 ;
        21:  q   <=  32'b00111111000001010111110011000111 ;
        22:  q   <=  32'b00111110111101001101110110110100 ;
        23:  q   <=  32'b00111110110111100010011000000010 ;
        24:  q   <=  32'b00111110110001101110000011101100 ;
        25:  q   <=  32'b00111110101011110001110101000011 ;
        26:  q   <=  32'b00111110100101101110101000100110 ;
        27:  q   <=  32'b00111110011111001010110111111000 ;
        28:  q   <=  32'b00111110010010101110011011010010 ;
        29:  q   <=  32'b00111110000110001001111010001001 ;
        30:  q   <=  32'b00111101110010111110101000111010 ;
        31:  q   <=  32'b00111101010011000010101100110011 ;
        32:  q   <=  32'b00100100100011010011000100110001 ;
        33:  q   <=  32'b10111101010011000010101100110011 ;
        34:  q   <=  32'b10111101110010111110101000111010 ;
        35:  q   <=  32'b10111110000110001001111010001001 ;
        36:  q   <=  32'b10111110010010101110011011010010 ;
        37:  q   <=  32'b10111110011111001010110111111000 ;
        38:  q   <=  32'b10111110100101101110101000100110 ;
        39:  q   <=  32'b10111110101011110001110101000011 ;
        40:  q   <=  32'b10111110110001101110000011101100 ;
        41:  q   <=  32'b10111110110111100010011000000010 ;
        42:  q   <=  32'b10111110111101001101110110110100 ;
        43:  q   <=  32'b10111111000001010111110011000111 ;
        44:  q   <=  32'b10111111000100000011010110111110 ;
        45:  q   <=  32'b10111111000110101001001011101101 ;
        46:  q   <=  32'b10111111001001001000110110111010 ;
        47:  q   <=  32'b10111111001011100001111111001100 ;
        48:  q   <=  32'b10111111001101110100001100001100 ;
        49:  q   <=  32'b10111111001111111111000110101001 ;
        50:  q   <=  32'b10111111010010000010011000011011 ;
        51:  q   <=  32'b10111111010011111101101100101011 ;
        52:  q   <=  32'b10111111010101110000101111110000 ;
        53:  q   <=  32'b10111111010111011011001111010111 ;
        54:  q   <=  32'b10111111011000111100111010100011 ;
        55:  q   <=  32'b10111111011010010101100001110010 ;
        56:  q   <=  32'b10111111011011100100110110111101 ;
        57:  q   <=  32'b10111111011100101010101101011101 ;
        58:  q   <=  32'b10111111011101100110111010001010 ;
        59:  q   <=  32'b10111111011110011001010011100000 ;
        60:  q   <=  32'b10111111011111000001110001011100 ;
        61:  q   <=  32'b10111111011111100000001101100011 ;
        62:  q   <=  32'b10111111011111110100100010111111 ;
        63:  q   <=  32'b10111111011111111110101110100001 ;
        64:  q   <=  32'b00111111011111111010111010001000 ;
        65:  q   <=  32'b00111111011111010010010000000100 ;
        66:  q   <=  32'b00111111011110000001010101110010 ;
        67:  q   <=  32'b00111111011100001000111110110010 ;
        68:  q   <=  32'b00111111011001101010010111100101 ;
        69:  q   <=  32'b00111111010110100111000101000101 ;
        70:  q   <=  32'b00111111010011000001000011100000 ;
        71:  q   <=  32'b00111111001110111010100101001001 ;
        72:  q   <=  32'b00111111001010010110010000111110 ;
        73:  q   <=  32'b00111111000101010111000000111001 ;
        74:  q   <=  32'b00111110111111111111111111111111 ;
        75:  q   <=  32'b00111110110100101001010000111001 ;
        76:  q   <=  32'b00111110101000110001000010101110 ;
        77:  q   <=  32'b00111110011000111101110010000111 ;
        78:  q   <=  32'b00111101111111101010011111101001 ;
        79:  q   <=  32'b00111100110011000011101101110011 ;
        80:  q   <=  32'b10111101100110010000110000010111 ;
        81:  q   <=  32'b10111110001100011101000011010011 ;
        82:  q   <=  32'b10111110100010101010101110011010 ;
        83:  q   <=  32'b10111110101110110000110111111010 ;
        84:  q   <=  32'b10111110111010011001010001110001 ;
        85:  q   <=  32'b10111111000010101110010001001111 ;
        86:  q   <=  32'b10111111000111111001110100000111 ;
        87:  q   <=  32'b10111111001100101011111110100101 ;
        88:  q   <=  32'b10111111010001000001101101111101 ;
        89:  q   <=  32'b10111111010100111000010001100010 ;
        90:  q   <=  32'b10111111011000001101001100100001 ;
        91:  q   <=  32'b10111111011010111110010111011101 ;
        92:  q   <=  32'b10111111011101001010000001101011 ;
        93:  q   <=  32'b10111111011110101110110010010101 ;
        94:  q   <=  32'b10111111011111101011101001010110 ;
        95:  q   <=  32'b10111111100000000000000000000000 ;
        96:  q   <=  32'b10111111011111101011101001010110 ;
        97:  q   <=  32'b10111111011110101110110010010101 ;
        98:  q   <=  32'b10111111011101001010000001101011 ;
        99:  q   <=  32'b10111111011010111110010111011101 ;
        100:  q   <=  32'b10111111011000001101001100100001 ;
        101:  q   <=  32'b10111111010100111000010001100010 ;
        102:  q   <=  32'b10111111010001000001101101111101 ;
        103:  q   <=  32'b10111111001100101011111110100101 ;
        104:  q   <=  32'b10111111000111111001110100000111 ;
        105:  q   <=  32'b10111111000010101110010001001111 ;
        106:  q   <=  32'b10111110111010011001010001110001 ;
        107:  q   <=  32'b10111110101110110000110111111010 ;
        108:  q   <=  32'b10111110100010101010101110011010 ;
        109:  q   <=  32'b10111110001100011101000011010011 ;
        110:  q   <=  32'b10111101100110010000110000010111 ;
        111:  q   <=  32'b00111100110011000011101101110011 ;
        112:  q   <=  32'b00111101111111101010011111101001 ;
        113:  q   <=  32'b00111110011000111101110010000111 ;
        114:  q   <=  32'b00111110101000110001000010101110 ;
        115:  q   <=  32'b00111110110100101001010000111001 ;
        116:  q   <=  32'b00111111000000000000000000000000 ;
        117:  q   <=  32'b00111111000101010111000000111001 ;
        118:  q   <=  32'b00111111001010010110010000111110 ;
        119:  q   <=  32'b00111111001110111010100101001001 ;
        120:  q   <=  32'b00111111010011000001000011100000 ;
        121:  q   <=  32'b00111111010110100111000101000101 ;
        122:  q   <=  32'b00111111011001101010010111100101 ;
        123:  q   <=  32'b00111111011100001000111110110010 ;
        124:  q   <=  32'b00111111011110000001010101110010 ;
        125:  q   <=  32'b00111111011111010010010000000100 ;
        126:  q   <=  32'b00111111011111111010111010001000 ;
        127:  q   <=  32'b00111111011111110100100010111111 ;
        128:  q   <=  32'b00111111011110011001010011100000 ;
        129:  q   <=  32'b00111111011011100100110110111101 ;
        130:  q   <=  32'b00111111010111011011001111010111 ;
        131:  q   <=  32'b00111111010010000010011000011011 ;
        132:  q   <=  32'b00111111001011100001111111001100 ;
        133:  q   <=  32'b00111111000100000011010110111110 ;
        134:  q   <=  32'b00111110110111100010011000000010 ;
        135:  q   <=  32'b00111110100101101110101000100110 ;
        136:  q   <=  32'b00111110000110001001111010001001 ;
        137:  q   <=  32'b00100100100011010011000100110001 ;
        138:  q   <=  32'b10111110000110001001111010001001 ;
        139:  q   <=  32'b10111110100101101110101000100110 ;
        140:  q   <=  32'b10111110110111100010011000000010 ;
        141:  q   <=  32'b10111111000100000011010110111110 ;
        142:  q   <=  32'b10111111001011100001111111001100 ;
        143:  q   <=  32'b10111111010010000010011000011011 ;
        144:  q   <=  32'b10111111010111011011001111010111 ;
        145:  q   <=  32'b10111111011011100100110110111101 ;
        146:  q   <=  32'b10111111011110011001010011100000 ;
        147:  q   <=  32'b10111111011111110100100010111111 ;
        148:  q   <=  32'b10111111011111110100100010111111 ;
        149:  q   <=  32'b10111111011110011001010011100000 ;
        150:  q   <=  32'b10111111011011100100110110111101 ;
        151:  q   <=  32'b10111111010111011011001111010111 ;
        152:  q   <=  32'b10111111010010000010011000011011 ;
        153:  q   <=  32'b10111111001011100001111111001100 ;
        154:  q   <=  32'b10111111000100000011010110111110 ;
        155:  q   <=  32'b10111110110111100010011000000010 ;
        156:  q   <=  32'b10111110100101101110101000100110 ;
        157:  q   <=  32'b10111110000110001001111010001001 ;
        158:  q   <=  32'b10100101010100111100100111001010 ;
        159:  q   <=  32'b00111110000110001001111010001001 ;
        160:  q   <=  32'b00111110100101101110101000100110 ;
        161:  q   <=  32'b00111110110111100010011000000010 ;
        162:  q   <=  32'b00111111000100000011010110111110 ;
        163:  q   <=  32'b00111111001011100001111111001100 ;
        164:  q   <=  32'b00111111010010000010011000011011 ;
        165:  q   <=  32'b00111111010111011011001111010111 ;
        166:  q   <=  32'b00111111011011100100110110111101 ;
        167:  q   <=  32'b00111111011110011001010011100000 ;
        168:  q   <=  32'b00111111011111110100100010111111 ;
        169:  q   <=  32'b00111111011111110100100010111111 ;
        170:  q   <=  32'b00111111011110011001010011100000 ;
        171:  q   <=  32'b00111111011011100100110110111101 ;
        172:  q   <=  32'b00111111010111011011001111010111 ;
        173:  q   <=  32'b00111111010010000010011000011011 ;
        174:  q   <=  32'b00111111001011100001111111001100 ;
        175:  q   <=  32'b00111111000100000011010110111110 ;
        176:  q   <=  32'b00111110110111100010011000000010 ;
        177:  q   <=  32'b00111110100101101110101000100110 ;
        178:  q   <=  32'b00111110000110001001111010001001 ;
        179:  q   <=  32'b00100101101100000111110101111101 ;
        180:  q   <=  32'b10111110000110001001111010001001 ;
        181:  q   <=  32'b10111110100101101110101000100110 ;
        182:  q   <=  32'b10111110110111100010011000000010 ;
        183:  q   <=  32'b10111111000100000011010110111110 ;
        184:  q   <=  32'b10111111001011100001111111001100 ;
        185:  q   <=  32'b10111111010010000010011000011011 ;
        186:  q   <=  32'b10111111010111011011001111010111 ;
        187:  q   <=  32'b10111111011011100100110110111101 ;
        188:  q   <=  32'b10111111011110011001010011100000 ;
        189:  q   <=  32'b10111111011111110100100010111111 ;
        190:  q   <=  32'b00111111011111101011101001010110 ;
        191:  q   <=  32'b00111111011101001010000001101011 ;
        192:  q   <=  32'b00111111011000001101001100100001 ;
        193:  q   <=  32'b00111111010001000001101101111101 ;
        194:  q   <=  32'b00111111000111111001110100000111 ;
        195:  q   <=  32'b00111110111010011001010001110001 ;
        196:  q   <=  32'b00111110100010101010101110011010 ;
        197:  q   <=  32'b00111101100110010000110000010111 ;
        198:  q   <=  32'b10111101111111101010011111101001 ;
        199:  q   <=  32'b10111110101000110001000010101110 ;
        200:  q   <=  32'b10111111000000000000000000000000 ;
        201:  q   <=  32'b10111111001010010110010000111110 ;
        202:  q   <=  32'b10111111010011000001000011100000 ;
        203:  q   <=  32'b10111111011001101010010111100101 ;
        204:  q   <=  32'b10111111011110000001010101110010 ;
        205:  q   <=  32'b10111111011111111010111010001000 ;
        206:  q   <=  32'b10111111011111010010010000000100 ;
        207:  q   <=  32'b10111111011100001000111110110010 ;
        208:  q   <=  32'b10111111010110100111000101000101 ;
        209:  q   <=  32'b10111111001110111010100101001001 ;
        210:  q   <=  32'b10111111000101010111000000111001 ;
        211:  q   <=  32'b10111110110100101001010000111001 ;
        212:  q   <=  32'b10111110011000111101110010000111 ;
        213:  q   <=  32'b10111100110011000011101101110011 ;
        214:  q   <=  32'b00111110001100011101000011010011 ;
        215:  q   <=  32'b00111110101110110000110111111010 ;
        216:  q   <=  32'b00111111000010101110010001001111 ;
        217:  q   <=  32'b00111111001100101011111110100101 ;
        218:  q   <=  32'b00111111010100111000010001100010 ;
        219:  q   <=  32'b00111111011010111110010111011101 ;
        220:  q   <=  32'b00111111011110101110110010010101 ;
        221:  q   <=  32'b00111111100000000000000000000000 ;
        222:  q   <=  32'b00111111011110101110110010010101 ;
        223:  q   <=  32'b00111111011010111110010111011101 ;
        224:  q   <=  32'b00111111010100111000010001100010 ;
        225:  q   <=  32'b00111111001100101011111110100101 ;
        226:  q   <=  32'b00111111000010101110010001001111 ;
        227:  q   <=  32'b00111110101110110000110111111010 ;
        228:  q   <=  32'b00111110001100011101000011010011 ;
        229:  q   <=  32'b10111100110011000011101101110011 ;
        230:  q   <=  32'b10111110011000111101110010000111 ;
        231:  q   <=  32'b10111110110100101001010000111001 ;
        232:  q   <=  32'b10111111000101010111000000111001 ;
        233:  q   <=  32'b10111111001110111010100101001001 ;
        234:  q   <=  32'b10111111010110100111000101000101 ;
        235:  q   <=  32'b10111111011100001000111110110010 ;
        236:  q   <=  32'b10111111011111010010010000000100 ;
        237:  q   <=  32'b10111111011111111010111010001000 ;
        238:  q   <=  32'b10111111011110000001010101110010 ;
        239:  q   <=  32'b10111111011001101010010111100101 ;
        240:  q   <=  32'b10111111010011000001000011100000 ;
        241:  q   <=  32'b10111111001010010110010000111110 ;
        242:  q   <=  32'b10111110111111111111111111111111 ;
        243:  q   <=  32'b10111110101000110001000010101110 ;
        244:  q   <=  32'b10111101111111101010011111101001 ;
        245:  q   <=  32'b00111101100110010000110000010111 ;
        246:  q   <=  32'b00111110100010101010101110011010 ;
        247:  q   <=  32'b00111110111010011001010001110001 ;
        248:  q   <=  32'b00111111000111111001110100000111 ;
        249:  q   <=  32'b00111111010001000001101101111101 ;
        250:  q   <=  32'b00111111011000001101001100100001 ;
        251:  q   <=  32'b00111111011101001010000001101011 ;
        252:  q   <=  32'b00111111011111101011101001010110 ;
        253:  q   <=  32'b00111111011111100000001101100011 ;
        254:  q   <=  32'b00111111011011100100110110111101 ;
        255:  q   <=  32'b00111111010011111101101100101011 ;
        256:  q   <=  32'b00111111001001001000110110111010 ;
        257:  q   <=  32'b00111110110111100010011000000010 ;
        258:  q   <=  32'b00111110010010101110011011010010 ;
        259:  q   <=  32'b10111101010011000010101100110011 ;
        260:  q   <=  32'b10111110100101101110101000100110 ;
        261:  q   <=  32'b10111111000001010111110011000111 ;
        262:  q   <=  32'b10111111001101110100001100001100 ;
        263:  q   <=  32'b10111111010111011011001111010111 ;
        264:  q   <=  32'b10111111011101100110111010001010 ;
        265:  q   <=  32'b10111111011111111110101110100001 ;
        266:  q   <=  32'b10111111011110011001010011100000 ;
        267:  q   <=  32'b10111111011000111100111010100011 ;
        268:  q   <=  32'b10111111001111111111000110101001 ;
        269:  q   <=  32'b10111111000100000011010110111110 ;
        270:  q   <=  32'b10111110101011110001110101000011 ;
        271:  q   <=  32'b10111101110010111110101000111010 ;
        272:  q   <=  32'b00111110000110001001111010001001 ;
        273:  q   <=  32'b00111110110001101110000011101100 ;
        274:  q   <=  32'b00111111000110101001001011101101 ;
        275:  q   <=  32'b00111111010010000010011000011011 ;
        276:  q   <=  32'b00111111011010010101100001110010 ;
        277:  q   <=  32'b00111111011111000001110001011100 ;
        278:  q   <=  32'b00111111011111110100100010111111 ;
        279:  q   <=  32'b00111111011100101010101101011101 ;
        280:  q   <=  32'b00111111010101110000101111110000 ;
        281:  q   <=  32'b00111111001011100001111111001100 ;
        282:  q   <=  32'b00111110111101001101110110110100 ;
        283:  q   <=  32'b00111110011111001010110111111000 ;
        284:  q   <=  32'b00100101101100000111110101111101 ;
        285:  q   <=  32'b10111110011111001010110111111000 ;
        286:  q   <=  32'b10111110111101001101110110110100 ;
        287:  q   <=  32'b10111111001011100001111111001100 ;
        288:  q   <=  32'b10111111010101110000101111110000 ;
        289:  q   <=  32'b10111111011100101010101101011101 ;
        290:  q   <=  32'b10111111011111110100100010111111 ;
        291:  q   <=  32'b10111111011111000001110001011100 ;
        292:  q   <=  32'b10111111011010010101100001110010 ;
        293:  q   <=  32'b10111111010010000010011000011011 ;
        294:  q   <=  32'b10111111000110101001001011101101 ;
        295:  q   <=  32'b10111110110001101110000011101100 ;
        296:  q   <=  32'b10111110000110001001111010001001 ;
        297:  q   <=  32'b00111101110010111110101000111010 ;
        298:  q   <=  32'b00111110101011110001110101000011 ;
        299:  q   <=  32'b00111111000100000011010110111110 ;
        300:  q   <=  32'b00111111001111111111000110101001 ;
        301:  q   <=  32'b00111111011000111100111010100011 ;
        302:  q   <=  32'b00111111011110011001010011100000 ;
        303:  q   <=  32'b00111111011111111110101110100001 ;
        304:  q   <=  32'b00111111011101100110111010001010 ;
        305:  q   <=  32'b00111111010111011011001111010111 ;
        306:  q   <=  32'b00111111001101110100001100001100 ;
        307:  q   <=  32'b00111111000001010111110011000111 ;
        308:  q   <=  32'b00111110100101101110101000100110 ;
        309:  q   <=  32'b00111101010011000010101100110011 ;
        310:  q   <=  32'b10111110010010101110011011010010 ;
        311:  q   <=  32'b10111110110111100010011000000010 ;
        312:  q   <=  32'b10111111001001001000110110111010 ;
        313:  q   <=  32'b10111111010011111101101100101011 ;
        314:  q   <=  32'b10111111011011100100110110111101 ;
        315:  q   <=  32'b10111111011111100000001101100011 ;
        316:  q   <=  32'b00111111011111010010010000000100 ;
        317:  q   <=  32'b00111111011001101010010111100101 ;
        318:  q   <=  32'b00111111001110111010100101001001 ;
        319:  q   <=  32'b00111110111111111111111111111111 ;
        320:  q   <=  32'b00111110011000111101110010000111 ;
        321:  q   <=  32'b10111101100110010000110000010111 ;
        322:  q   <=  32'b10111110101110110000110111111010 ;
        323:  q   <=  32'b10111111000111111001110100000111 ;
        324:  q   <=  32'b10111111010100111000010001100010 ;
        325:  q   <=  32'b10111111011101001010000001101011 ;
        326:  q   <=  32'b10111111100000000000000000000000 ;
        327:  q   <=  32'b10111111011101001010000001101011 ;
        328:  q   <=  32'b10111111010100111000010001100010 ;
        329:  q   <=  32'b10111111000111111001110100000111 ;
        330:  q   <=  32'b10111110101110110000110111111010 ;
        331:  q   <=  32'b10111101100110010000110000010111 ;
        332:  q   <=  32'b00111110011000111101110010000111 ;
        333:  q   <=  32'b00111111000000000000000000000000 ;
        334:  q   <=  32'b00111111001110111010100101001001 ;
        335:  q   <=  32'b00111111011001101010010111100101 ;
        336:  q   <=  32'b00111111011111010010010000000100 ;
        337:  q   <=  32'b00111111011111010010010000000100 ;
        338:  q   <=  32'b00111111011001101010010111100101 ;
        339:  q   <=  32'b00111111001110111010100101001001 ;
        340:  q   <=  32'b00111110111111111111111111111111 ;
        341:  q   <=  32'b00111110011000111101110010000111 ;
        342:  q   <=  32'b10111101100110010000110000010111 ;
        343:  q   <=  32'b10111110101110110000110111111010 ;
        344:  q   <=  32'b10111111000111111001110100000111 ;
        345:  q   <=  32'b10111111010100111000010001100010 ;
        346:  q   <=  32'b10111111011101001010000001101011 ;
        347:  q   <=  32'b10111111100000000000000000000000 ;
        348:  q   <=  32'b10111111011101001010000001101011 ;
        349:  q   <=  32'b10111111010100111000010001100010 ;
        350:  q   <=  32'b10111111000111111001110100000111 ;
        351:  q   <=  32'b10111110101110110000110111111010 ;
        352:  q   <=  32'b10111101100110010000110000010111 ;
        353:  q   <=  32'b00111110011000111101110010000111 ;
        354:  q   <=  32'b00111111000000000000000000000000 ;
        355:  q   <=  32'b00111111001110111010100101001001 ;
        356:  q   <=  32'b00111111011001101010010111100101 ;
        357:  q   <=  32'b00111111011111010010010000000100 ;
        358:  q   <=  32'b00111111011111010010010000000100 ;
        359:  q   <=  32'b00111111011001101010010111100101 ;
        360:  q   <=  32'b00111111001110111010100101001001 ;
        361:  q   <=  32'b00111110111111111111111111111111 ;
        362:  q   <=  32'b00111110011000111101110010000111 ;
        363:  q   <=  32'b10111101100110010000110000010111 ;
        364:  q   <=  32'b10111110101110110000110111111010 ;
        365:  q   <=  32'b10111111000111111001110100000111 ;
        366:  q   <=  32'b10111111010100111000010001100010 ;
        367:  q   <=  32'b10111111011101001010000001101011 ;
        368:  q   <=  32'b10111111100000000000000000000000 ;
        369:  q   <=  32'b10111111011101001010000001101011 ;
        370:  q   <=  32'b10111111010100111000010001100010 ;
        371:  q   <=  32'b10111111000111111001110100000111 ;
        372:  q   <=  32'b10111110101110110000110111111010 ;
        373:  q   <=  32'b10111101100110010000110000010111 ;
        374:  q   <=  32'b00111110011000111101110010000111 ;
        375:  q   <=  32'b00111110111111111111111111111111 ;
        376:  q   <=  32'b00111111001110111010100101001001 ;
        377:  q   <=  32'b00111111011001101010010111100101 ;
        378:  q   <=  32'b00111111011111010010010000000100 ;
        379:  q   <=  32'b00111111011111000001110001011100 ;
        380:  q   <=  32'b00111111010111011011001111010111 ;
        381:  q   <=  32'b00111111001001001000110110111010 ;
        382:  q   <=  32'b00111110101011110001110101000011 ;
        383:  q   <=  32'b00100100100011010011000100110001 ;
        384:  q   <=  32'b10111110101011110001110101000011 ;
        385:  q   <=  32'b10111111001001001000110110111010 ;
        386:  q   <=  32'b10111111010111011011001111010111 ;
        387:  q   <=  32'b10111111011111000001110001011100 ;
        388:  q   <=  32'b10111111011111000001110001011100 ;
        389:  q   <=  32'b10111111010111011011001111010111 ;
        390:  q   <=  32'b10111111001001001000110110111010 ;
        391:  q   <=  32'b10111110101011110001110101000011 ;
        392:  q   <=  32'b10100101010100111100100111001010 ;
        393:  q   <=  32'b00111110101011110001110101000011 ;
        394:  q   <=  32'b00111111001001001000110110111010 ;
        395:  q   <=  32'b00111111010111011011001111010111 ;
        396:  q   <=  32'b00111111011111000001110001011100 ;
        397:  q   <=  32'b00111111011111000001110001011100 ;
        398:  q   <=  32'b00111111010111011011001111010111 ;
        399:  q   <=  32'b00111111001001001000110110111010 ;
        400:  q   <=  32'b00111110101011110001110101000011 ;
        401:  q   <=  32'b00100101101100000111110101111101 ;
        402:  q   <=  32'b10111110101011110001110101000011 ;
        403:  q   <=  32'b10111111001001001000110110111010 ;
        404:  q   <=  32'b10111111010111011011001111010111 ;
        405:  q   <=  32'b10111111011111000001110001011100 ;
        406:  q   <=  32'b10111111011111000001110001011100 ;
        407:  q   <=  32'b10111111010111011011001111010111 ;
        408:  q   <=  32'b10111111001001001000110110111010 ;
        409:  q   <=  32'b10111110101011110001110101000011 ;
        410:  q   <=  32'b10100101111101110001011000010110 ;
        411:  q   <=  32'b00111110101011110001110101000011 ;
        412:  q   <=  32'b00111111001001001000110110111010 ;
        413:  q   <=  32'b00111111010111011011001111010111 ;
        414:  q   <=  32'b00111111011111000001110001011100 ;
        415:  q   <=  32'b00111111011111000001110001011100 ;
        416:  q   <=  32'b00111111010111011011001111010111 ;
        417:  q   <=  32'b00111111001001001000110110111010 ;
        418:  q   <=  32'b00111110101011110001110101000011 ;
        419:  q   <=  32'b00100110000111101101011101010111 ;
        420:  q   <=  32'b10111110101011110001110101000011 ;
        421:  q   <=  32'b10111111001001001000110110111010 ;
        422:  q   <=  32'b10111111010111011011001111010111 ;
        423:  q   <=  32'b10111111011111000001110001011100 ;
        424:  q   <=  32'b10111111011111000001110001011100 ;
        425:  q   <=  32'b10111111010111011011001111010111 ;
        426:  q   <=  32'b10111111001001001000110110111010 ;
        427:  q   <=  32'b10111110101011110001110101000011 ;
        428:  q   <=  32'b10100111001100001000100011101001 ;
        429:  q   <=  32'b00111110101011110001110101000011 ;
        430:  q   <=  32'b00111111001001001000110110111010 ;
        431:  q   <=  32'b00111111010111011011001111010111 ;
        432:  q   <=  32'b00111111011111000001110001011100 ;
        433:  q   <=  32'b00111111011111000001110001011100 ;
        434:  q   <=  32'b00111111010111011011001111010111 ;
        435:  q   <=  32'b00111111001001001000110110111010 ;
        436:  q   <=  32'b00111110101011110001110101000011 ;
        437:  q   <=  32'b10100110100011010100100000000111 ;
        438:  q   <=  32'b10111110101011110001110101000011 ;
        439:  q   <=  32'b10111111001001001000110110111010 ;
        440:  q   <=  32'b10111111010111011011001111010111 ;
        441:  q   <=  32'b10111111011111000001110001011100 ;
        442:  q   <=  32'b00111111011110101110110010010101 ;
        443:  q   <=  32'b00111111010100111000010001100010 ;
        444:  q   <=  32'b00111111000010101110010001001111 ;
        445:  q   <=  32'b00111110001100011101000011010011 ;
        446:  q   <=  32'b10111110011000111101110010000111 ;
        447:  q   <=  32'b10111111000101010111000000111001 ;
        448:  q   <=  32'b10111111010110100111000101000101 ;
        449:  q   <=  32'b10111111011111010010010000000100 ;
        450:  q   <=  32'b10111111011110000001010101110010 ;
        451:  q   <=  32'b10111111010011000001000011100000 ;
        452:  q   <=  32'b10111110111111111111111111111111 ;
        453:  q   <=  32'b10111101111111101010011111101001 ;
        454:  q   <=  32'b00111110100010101010101110011010 ;
        455:  q   <=  32'b00111111000111111001110100000111 ;
        456:  q   <=  32'b00111111011000001101001100100001 ;
        457:  q   <=  32'b00111111011111101011101001010110 ;
        458:  q   <=  32'b00111111011101001010000001101011 ;
        459:  q   <=  32'b00111111010001000001101101111101 ;
        460:  q   <=  32'b00111110111010011001010001110001 ;
        461:  q   <=  32'b00111101100110010000110000010111 ;
        462:  q   <=  32'b10111110101000110001000010101110 ;
        463:  q   <=  32'b10111111001010010110010000111110 ;
        464:  q   <=  32'b10111111011001101010010111100101 ;
        465:  q   <=  32'b10111111011111111010111010001000 ;
        466:  q   <=  32'b10111111011100001000111110110010 ;
        467:  q   <=  32'b10111111001110111010100101001001 ;
        468:  q   <=  32'b10111110110100101001010000111001 ;
        469:  q   <=  32'b10111100110011000011101101110011 ;
        470:  q   <=  32'b00111110101110110000110111111010 ;
        471:  q   <=  32'b00111111001100101011111110100101 ;
        472:  q   <=  32'b00111111011010111110010111011101 ;
        473:  q   <=  32'b00111111100000000000000000000000 ;
        474:  q   <=  32'b00111111011010111110010111011101 ;
        475:  q   <=  32'b00111111001100101011111110100101 ;
        476:  q   <=  32'b00111110101110110000110111111010 ;
        477:  q   <=  32'b10111100110011000011101101110011 ;
        478:  q   <=  32'b10111110110100101001010000111001 ;
        479:  q   <=  32'b10111111001110111010100101001001 ;
        480:  q   <=  32'b10111111011100001000111110110010 ;
        481:  q   <=  32'b10111111011111111010111010001000 ;
        482:  q   <=  32'b10111111011001101010010111100101 ;
        483:  q   <=  32'b10111111001010010110010000111110 ;
        484:  q   <=  32'b10111110101000110001000010101110 ;
        485:  q   <=  32'b00111101100110010000110000010111 ;
        486:  q   <=  32'b00111110111010011001010001110001 ;
        487:  q   <=  32'b00111111010001000001101101111101 ;
        488:  q   <=  32'b00111111011101001010000001101011 ;
        489:  q   <=  32'b00111111011111101011101001010110 ;
        490:  q   <=  32'b00111111011000001101001100100001 ;
        491:  q   <=  32'b00111111000111111001110100000111 ;
        492:  q   <=  32'b00111110100010101010101110011010 ;
        493:  q   <=  32'b10111101111111101010011111101001 ;
        494:  q   <=  32'b10111111000000000000000000000000 ;
        495:  q   <=  32'b10111111010011000001000011100000 ;
        496:  q   <=  32'b10111111011110000001010101110010 ;
        497:  q   <=  32'b10111111011111010010010000000100 ;
        498:  q   <=  32'b10111111010110100111000101000101 ;
        499:  q   <=  32'b10111111000101010111000000111001 ;
        500:  q   <=  32'b10111110011000111101110010000111 ;
        501:  q   <=  32'b00111110001100011101000011010011 ;
        502:  q   <=  32'b00111111000010101110010001001111 ;
        503:  q   <=  32'b00111111010100111000010001100010 ;
        504:  q   <=  32'b00111111011110101110110010010101 ;
        505:  q   <=  32'b00111111011110011001010011100000 ;
        506:  q   <=  32'b00111111010010000010011000011011 ;
        507:  q   <=  32'b00111110110111100010011000000010 ;
        508:  q   <=  32'b00100100100011010011000100110001 ;
        509:  q   <=  32'b10111110110111100010011000000010 ;
        510:  q   <=  32'b10111111010010000010011000011011 ;
        511:  q   <=  32'b10111111011110011001010011100000 ;
        512:  q   <=  32'b10111111011110011001010011100000 ;
        513:  q   <=  32'b10111111010010000010011000011011 ;
        514:  q   <=  32'b10111110110111100010011000000010 ;
        515:  q   <=  32'b10100101010100111100100111001010 ;
        516:  q   <=  32'b00111110110111100010011000000010 ;
        517:  q   <=  32'b00111111010010000010011000011011 ;
        518:  q   <=  32'b00111111011110011001010011100000 ;
        519:  q   <=  32'b00111111011110011001010011100000 ;
        520:  q   <=  32'b00111111010010000010011000011011 ;
        521:  q   <=  32'b00111110110111100010011000000010 ;
        522:  q   <=  32'b00100101101100000111110101111101 ;
        523:  q   <=  32'b10111110110111100010011000000010 ;
        524:  q   <=  32'b10111111010010000010011000011011 ;
        525:  q   <=  32'b10111111011110011001010011100000 ;
        526:  q   <=  32'b10111111011110011001010011100000 ;
        527:  q   <=  32'b10111111010010000010011000011011 ;
        528:  q   <=  32'b10111110110111100010011000000010 ;
        529:  q   <=  32'b10100101111101110001011000010110 ;
        530:  q   <=  32'b00111110110111100010011000000010 ;
        531:  q   <=  32'b00111111010010000010011000011011 ;
        532:  q   <=  32'b00111111011110011001010011100000 ;
        533:  q   <=  32'b00111111011110011001010011100000 ;
        534:  q   <=  32'b00111111010010000010011000011011 ;
        535:  q   <=  32'b00111110110111100010011000000010 ;
        536:  q   <=  32'b00100110000111101101011101010111 ;
        537:  q   <=  32'b10111110110111100010011000000010 ;
        538:  q   <=  32'b10111111010010000010011000011011 ;
        539:  q   <=  32'b10111111011110011001010011100000 ;
        540:  q   <=  32'b10111111011110011001010011100000 ;
        541:  q   <=  32'b10111111010010000010011000011011 ;
        542:  q   <=  32'b10111110110111100010011000000010 ;
        543:  q   <=  32'b10100111001100001000100011101001 ;
        544:  q   <=  32'b00111110110111100010011000000010 ;
        545:  q   <=  32'b00111111010010000010011000011011 ;
        546:  q   <=  32'b00111111011110011001010011100000 ;
        547:  q   <=  32'b00111111011110011001010011100000 ;
        548:  q   <=  32'b00111111010010000010011000011011 ;
        549:  q   <=  32'b00111110110111100010011000000010 ;
        550:  q   <=  32'b10100110100011010100100000000111 ;
        551:  q   <=  32'b10111110110111100010011000000010 ;
        552:  q   <=  32'b10111111010010000010011000011011 ;
        553:  q   <=  32'b10111111011110011001010011100000 ;
        554:  q   <=  32'b10111111011110011001010011100000 ;
        555:  q   <=  32'b10111111010010000010011000011011 ;
        556:  q   <=  32'b10111110110111100010011000000010 ;
        557:  q   <=  32'b10100111010000100010111100001111 ;
        558:  q   <=  32'b00111110110111100010011000000010 ;
        559:  q   <=  32'b00111111010010000010011000011011 ;
        560:  q   <=  32'b00111111011110011001010011100000 ;
        561:  q   <=  32'b00111111011110011001010011100000 ;
        562:  q   <=  32'b00111111010010000010011000011011 ;
        563:  q   <=  32'b00111110110111100010011000000010 ;
        564:  q   <=  32'b10100110010100111111011101110110 ;
        565:  q   <=  32'b10111110110111100010011000000010 ;
        566:  q   <=  32'b10111111010010000010011000011011 ;
        567:  q   <=  32'b10111111011110011001010011100000 ;
        568:  q   <=  32'b00111111011110000001010101110010 ;
        569:  q   <=  32'b00111111001110111010100101001001 ;
        570:  q   <=  32'b00111110101000110001000010101110 ;
        571:  q   <=  32'b10111110001100011101000011010011 ;
        572:  q   <=  32'b10111111000111111001110100000111 ;
        573:  q   <=  32'b10111111011010111110010111011101 ;
        574:  q   <=  32'b10111111011111101011101001010110 ;
        575:  q   <=  32'b10111111010100111000010001100010 ;
        576:  q   <=  32'b10111110111010011001010001110001 ;
        577:  q   <=  32'b00111100110011000011101101110011 ;
        578:  q   <=  32'b00111111000000000000000000000000 ;
        579:  q   <=  32'b00111111010110100111000101000101 ;
        580:  q   <=  32'b00111111011111111010111010001000 ;
        581:  q   <=  32'b00111111011001101010010111100101 ;
        582:  q   <=  32'b00111111000101010111000000111001 ;
        583:  q   <=  32'b00111101111111101010011111101001 ;
        584:  q   <=  32'b10111110101110110000110111111010 ;
        585:  q   <=  32'b10111111010001000001101101111101 ;
        586:  q   <=  32'b10111111011110101110110010010101 ;
        587:  q   <=  32'b10111111011101001010000001101011 ;
        588:  q   <=  32'b10111111001100101011111110100101 ;
        589:  q   <=  32'b10111110100010101010101110011010 ;
        590:  q   <=  32'b00111110011000111101110010000111 ;
        591:  q   <=  32'b00111111001010010110010000111110 ;
        592:  q   <=  32'b00111111011100001000111110110010 ;
        593:  q   <=  32'b00111111011111010010010000000100 ;
        594:  q   <=  32'b00111111010011000001000011100000 ;
        595:  q   <=  32'b00111110110100101001010000111001 ;
        596:  q   <=  32'b10111101100110010000110000010111 ;
        597:  q   <=  32'b10111111000010101110010001001111 ;
        598:  q   <=  32'b10111111011000001101001100100001 ;
        599:  q   <=  32'b10111111100000000000000000000000 ;
        600:  q   <=  32'b10111111011000001101001100100001 ;
        601:  q   <=  32'b10111111000010101110010001001111 ;
        602:  q   <=  32'b10111101100110010000110000010111 ;
        603:  q   <=  32'b00111110110100101001010000111001 ;
        604:  q   <=  32'b00111111010011000001000011100000 ;
        605:  q   <=  32'b00111111011111010010010000000100 ;
        606:  q   <=  32'b00111111011100001000111110110010 ;
        607:  q   <=  32'b00111111001010010110010000111110 ;
        608:  q   <=  32'b00111110011000111101110010000111 ;
        609:  q   <=  32'b10111110100010101010101110011010 ;
        610:  q   <=  32'b10111111001100101011111110100101 ;
        611:  q   <=  32'b10111111011101001010000001101011 ;
        612:  q   <=  32'b10111111011110101110110010010101 ;
        613:  q   <=  32'b10111111010001000001101101111101 ;
        614:  q   <=  32'b10111110101110110000110111111010 ;
        615:  q   <=  32'b00111101111111101010011111101001 ;
        616:  q   <=  32'b00111111000101010111000000111001 ;
        617:  q   <=  32'b00111111011001101010010111100101 ;
        618:  q   <=  32'b00111111011111111010111010001000 ;
        619:  q   <=  32'b00111111010110100111000101000101 ;
        620:  q   <=  32'b00111111000000000000000000000000 ;
        621:  q   <=  32'b00111100110011000011101101110011 ;
        622:  q   <=  32'b10111110111010011001010001110001 ;
        623:  q   <=  32'b10111111010100111000010001100010 ;
        624:  q   <=  32'b10111111011111101011101001010110 ;
        625:  q   <=  32'b10111111011010111110010111011101 ;
        626:  q   <=  32'b10111111000111111001110100000111 ;
        627:  q   <=  32'b10111110001100011101000011010011 ;
        628:  q   <=  32'b00111110101000110001000010101110 ;
        629:  q   <=  32'b00111111001110111010100101001001 ;
        630:  q   <=  32'b00111111011110000001010101110010 ;
        631:  q   <=  32'b00111111011101100110111010001010 ;
        632:  q   <=  32'b00111111001011100001111111001100 ;
        633:  q   <=  32'b00111110010010101110011011010010 ;
        634:  q   <=  32'b10111110101011110001110101000011 ;
        635:  q   <=  32'b10111111010010000010011000011011 ;
        636:  q   <=  32'b10111111011111100000001101100011 ;
        637:  q   <=  32'b10111111011010010101100001110010 ;
        638:  q   <=  32'b10111111000100000011010110111110 ;
        639:  q   <=  32'b10111101010011000010101100110011 ;
        640:  q   <=  32'b00111110111101001101110110110100 ;
        641:  q   <=  32'b00111111010111011011001111010111 ;
        642:  q   <=  32'b00111111011111111110101110100001 ;
        643:  q   <=  32'b00111111010101110000101111110000 ;
        644:  q   <=  32'b00111110110111100010011000000010 ;
        645:  q   <=  32'b10111101110010111110101000111010 ;
        646:  q   <=  32'b10111111000110101001001011101101 ;
        647:  q   <=  32'b10111111011011100100110110111101 ;
        648:  q   <=  32'b10111111011111000001110001011100 ;
        649:  q   <=  32'b10111111001111111111000110101001 ;
        650:  q   <=  32'b10111110100101101110101000100110 ;
        651:  q   <=  32'b00111110011111001010110111111000 ;
        652:  q   <=  32'b00111111001101110100001100001100 ;
        653:  q   <=  32'b00111111011110011001010011100000 ;
        654:  q   <=  32'b00111111011100101010101101011101 ;
        655:  q   <=  32'b00111111001001001000110110111010 ;
        656:  q   <=  32'b00111110000110001001111010001001 ;
        657:  q   <=  32'b10111110110001101110000011101100 ;
        658:  q   <=  32'b10111111010011111101101100101011 ;
        659:  q   <=  32'b10111111011111110100100010111111 ;
        660:  q   <=  32'b10111111011000111100111010100011 ;
        661:  q   <=  32'b10111111000001010111110011000111 ;
        662:  q   <=  32'b10100111001100001000100011101001 ;
        663:  q   <=  32'b00111111000001010111110011000111 ;
        664:  q   <=  32'b00111111011000111100111010100011 ;
        665:  q   <=  32'b00111111011111110100100010111111 ;
        666:  q   <=  32'b00111111010011111101101100101011 ;
        667:  q   <=  32'b00111110110001101110000011101100 ;
        668:  q   <=  32'b10111110000110001001111010001001 ;
        669:  q   <=  32'b10111111001001001000110110111010 ;
        670:  q   <=  32'b10111111011100101010101101011101 ;
        671:  q   <=  32'b10111111011110011001010011100000 ;
        672:  q   <=  32'b10111111001101110100001100001100 ;
        673:  q   <=  32'b10111110011111001010110111111000 ;
        674:  q   <=  32'b00111110100101101110101000100110 ;
        675:  q   <=  32'b00111111001111111111000110101001 ;
        676:  q   <=  32'b00111111011111000001110001011100 ;
        677:  q   <=  32'b00111111011011100100110110111101 ;
        678:  q   <=  32'b00111111000110101001001011101101 ;
        679:  q   <=  32'b00111101110010111110101000111010 ;
        680:  q   <=  32'b10111110110111100010011000000010 ;
        681:  q   <=  32'b10111111010101110000101111110000 ;
        682:  q   <=  32'b10111111011111111110101110100001 ;
        683:  q   <=  32'b10111111010111011011001111010111 ;
        684:  q   <=  32'b10111110111101001101110110110100 ;
        685:  q   <=  32'b00111101010011000010101100110011 ;
        686:  q   <=  32'b00111111000100000011010110111110 ;
        687:  q   <=  32'b00111111011010010101100001110010 ;
        688:  q   <=  32'b00111111011111100000001101100011 ;
        689:  q   <=  32'b00111111010010000010011000011011 ;
        690:  q   <=  32'b00111110101011110001110101000011 ;
        691:  q   <=  32'b10111110010010101110011011010010 ;
        692:  q   <=  32'b10111111001011100001111111001100 ;
        693:  q   <=  32'b10111111011101100110111010001010 ;
        694:  q   <=  32'b00111111011101001010000001101011 ;
        695:  q   <=  32'b00111111000111111001110100000111 ;
        696:  q   <=  32'b00111101100110010000110000010111 ;
        697:  q   <=  32'b10111111000000000000000000000000 ;
        698:  q   <=  32'b10111111011001101010010111100101 ;
        699:  q   <=  32'b10111111011111010010010000000100 ;
        700:  q   <=  32'b10111111001110111010100101001001 ;
        701:  q   <=  32'b10111110011000111101110010000111 ;
        702:  q   <=  32'b00111110101110110000110111111010 ;
        703:  q   <=  32'b00111111010100111000010001100010 ;
        704:  q   <=  32'b00111111100000000000000000000000 ;
        705:  q   <=  32'b00111111010100111000010001100010 ;
        706:  q   <=  32'b00111110101110110000110111111010 ;
        707:  q   <=  32'b10111110011000111101110010000111 ;
        708:  q   <=  32'b10111111001110111010100101001001 ;
        709:  q   <=  32'b10111111011111010010010000000100 ;
        710:  q   <=  32'b10111111011001101010010111100101 ;
        711:  q   <=  32'b10111110111111111111111111111111 ;
        712:  q   <=  32'b00111101100110010000110000010111 ;
        713:  q   <=  32'b00111111000111111001110100000111 ;
        714:  q   <=  32'b00111111011101001010000001101011 ;
        715:  q   <=  32'b00111111011101001010000001101011 ;
        716:  q   <=  32'b00111111000111111001110100000111 ;
        717:  q   <=  32'b00111101100110010000110000010111 ;
        718:  q   <=  32'b10111111000000000000000000000000 ;
        719:  q   <=  32'b10111111011001101010010111100101 ;
        720:  q   <=  32'b10111111011111010010010000000100 ;
        721:  q   <=  32'b10111111001110111010100101001001 ;
        722:  q   <=  32'b10111110011000111101110010000111 ;
        723:  q   <=  32'b00111110101110110000110111111010 ;
        724:  q   <=  32'b00111111010100111000010001100010 ;
        725:  q   <=  32'b00111111100000000000000000000000 ;
        726:  q   <=  32'b00111111010100111000010001100010 ;
        727:  q   <=  32'b00111110101110110000110111111010 ;
        728:  q   <=  32'b10111110011000111101110010000111 ;
        729:  q   <=  32'b10111111001110111010100101001001 ;
        730:  q   <=  32'b10111111011111010010010000000100 ;
        731:  q   <=  32'b10111111011001101010010111100101 ;
        732:  q   <=  32'b10111110111111111111111111111111 ;
        733:  q   <=  32'b00111101100110010000110000010111 ;
        734:  q   <=  32'b00111111000111111001110100000111 ;
        735:  q   <=  32'b00111111011101001010000001101011 ;
        736:  q   <=  32'b00111111011101001010000001101011 ;
        737:  q   <=  32'b00111111000111111001110100000111 ;
        738:  q   <=  32'b00111101100110010000110000010111 ;
        739:  q   <=  32'b10111111000000000000000000000000 ;
        740:  q   <=  32'b10111111011001101010010111100101 ;
        741:  q   <=  32'b10111111011111010010010000000100 ;
        742:  q   <=  32'b10111111001110111010100101001001 ;
        743:  q   <=  32'b10111110011000111101110010000111 ;
        744:  q   <=  32'b00111110101110110000110111111010 ;
        745:  q   <=  32'b00111111010100111000010001100010 ;
        746:  q   <=  32'b00111111100000000000000000000000 ;
        747:  q   <=  32'b00111111010100111000010001100010 ;
        748:  q   <=  32'b00111110101110110000110111111010 ;
        749:  q   <=  32'b10111110011000111101110010000111 ;
        750:  q   <=  32'b10111111001110111010100101001001 ;
        751:  q   <=  32'b10111111011111010010010000000100 ;
        752:  q   <=  32'b10111111011001101010010111100101 ;
        753:  q   <=  32'b10111111000000000000000000000000 ;
        754:  q   <=  32'b00111101100110010000110000010111 ;
        755:  q   <=  32'b00111111000111111001110100000111 ;
        756:  q   <=  32'b00111111011101001010000001101011 ;
        757:  q   <=  32'b00111111011100101010101101011101 ;
        758:  q   <=  32'b00111111000100000011010110111110 ;
        759:  q   <=  32'b10111101010011000010101100110011 ;
        760:  q   <=  32'b10111111001001001000110110111010 ;
        761:  q   <=  32'b10111111011110011001010011100000 ;
        762:  q   <=  32'b10111111011010010101100001110010 ;
        763:  q   <=  32'b10111110111101001101110110110100 ;
        764:  q   <=  32'b00111110000110001001111010001001 ;
        765:  q   <=  32'b00111111001101110100001100001100 ;
        766:  q   <=  32'b00111111011111100000001101100011 ;
        767:  q   <=  32'b00111111010111011011001111010111 ;
        768:  q   <=  32'b00111110110001101110000011101100 ;
        769:  q   <=  32'b10111110011111001010110111111000 ;
        770:  q   <=  32'b10111111010010000010011000011011 ;
        771:  q   <=  32'b10111111011111111110101110100001 ;
        772:  q   <=  32'b10111111010011111101101100101011 ;
        773:  q   <=  32'b10111110100101101110101000100110 ;
        774:  q   <=  32'b00111110101011110001110101000011 ;
        775:  q   <=  32'b00111111010101110000101111110000 ;
        776:  q   <=  32'b00111111011111110100100010111111 ;
        777:  q   <=  32'b00111111001111111111000110101001 ;
        778:  q   <=  32'b00111110010010101110011011010010 ;
        779:  q   <=  32'b10111110110111100010011000000010 ;
        780:  q   <=  32'b10111111011000111100111010100011 ;
        781:  q   <=  32'b10111111011111000001110001011100 ;
        782:  q   <=  32'b10111111001011100001111111001100 ;
        783:  q   <=  32'b10111101110010111110101000111010 ;
        784:  q   <=  32'b00111111000001010111110011000111 ;
        785:  q   <=  32'b00111111011011100100110110111101 ;
        786:  q   <=  32'b00111111011101100110111010001010 ;
        787:  q   <=  32'b00111111000110101001001011101101 ;
        788:  q   <=  32'b10100110100011010100100000000111 ;
        789:  q   <=  32'b10111111000110101001001011101101 ;
        790:  q   <=  32'b10111111011101100110111010001010 ;
        791:  q   <=  32'b10111111011011100100110110111101 ;
        792:  q   <=  32'b10111111000001010111110011000111 ;
        793:  q   <=  32'b00111101110010111110101000111010 ;
        794:  q   <=  32'b00111111001011100001111111001100 ;
        795:  q   <=  32'b00111111011111000001110001011100 ;
        796:  q   <=  32'b00111111011000111100111010100011 ;
        797:  q   <=  32'b00111110110111100010011000000010 ;
        798:  q   <=  32'b10111110010010101110011011010010 ;
        799:  q   <=  32'b10111111001111111111000110101001 ;
        800:  q   <=  32'b10111111011111110100100010111111 ;
        801:  q   <=  32'b10111111010101110000101111110000 ;
        802:  q   <=  32'b10111110101011110001110101000011 ;
        803:  q   <=  32'b00111110100101101110101000100110 ;
        804:  q   <=  32'b00111111010011111101101100101011 ;
        805:  q   <=  32'b00111111011111111110101110100001 ;
        806:  q   <=  32'b00111111010010000010011000011011 ;
        807:  q   <=  32'b00111110011111001010110111111000 ;
        808:  q   <=  32'b10111110110001101110000011101100 ;
        809:  q   <=  32'b10111111010111011011001111010111 ;
        810:  q   <=  32'b10111111011111100000001101100011 ;
        811:  q   <=  32'b10111111001101110100001100001100 ;
        812:  q   <=  32'b10111110000110001001111010001001 ;
        813:  q   <=  32'b00111110111101001101110110110100 ;
        814:  q   <=  32'b00111111011010010101100001110010 ;
        815:  q   <=  32'b00111111011110011001010011100000 ;
        816:  q   <=  32'b00111111001001001000110110111010 ;
        817:  q   <=  32'b00111101010011000010101100110011 ;
        818:  q   <=  32'b10111111000100000011010110111110 ;
        819:  q   <=  32'b10111111011100101010101101011101 ;
        820:  q   <=  32'b00111111011100001000111110110010 ;
        821:  q   <=  32'b00111110111111111111111111111111 ;
        822:  q   <=  32'b10111110001100011101000011010011 ;
        823:  q   <=  32'b10111111010001000001101101111101 ;
        824:  q   <=  32'b10111111100000000000000000000000 ;
        825:  q   <=  32'b10111111010001000001101101111101 ;
        826:  q   <=  32'b10111110001100011101000011010011 ;
        827:  q   <=  32'b00111111000000000000000000000000 ;
        828:  q   <=  32'b00111111011100001000111110110010 ;
        829:  q   <=  32'b00111111011100001000111110110010 ;
        830:  q   <=  32'b00111110111111111111111111111111 ;
        831:  q   <=  32'b10111110001100011101000011010011 ;
        832:  q   <=  32'b10111111010001000001101101111101 ;
        833:  q   <=  32'b10111111100000000000000000000000 ;
        834:  q   <=  32'b10111111010001000001101101111101 ;
        835:  q   <=  32'b10111110001100011101000011010011 ;
        836:  q   <=  32'b00111111000000000000000000000000 ;
        837:  q   <=  32'b00111111011100001000111110110010 ;
        838:  q   <=  32'b00111111011100001000111110110010 ;
        839:  q   <=  32'b00111110111111111111111111111111 ;
        840:  q   <=  32'b10111110001100011101000011010011 ;
        841:  q   <=  32'b10111111010001000001101101111101 ;
        842:  q   <=  32'b10111111100000000000000000000000 ;
        843:  q   <=  32'b10111111010001000001101101111101 ;
        844:  q   <=  32'b10111110001100011101000011010011 ;
        845:  q   <=  32'b00111110111111111111111111111111 ;
        846:  q   <=  32'b00111111011100001000111110110010 ;
        847:  q   <=  32'b00111111011100001000111110110010 ;
        848:  q   <=  32'b00111111000000000000000000000000 ;
        849:  q   <=  32'b10111110001100011101000011010011 ;
        850:  q   <=  32'b10111111010001000001101101111101 ;
        851:  q   <=  32'b10111111100000000000000000000000 ;
        852:  q   <=  32'b10111111010001000001101101111101 ;
        853:  q   <=  32'b10111110001100011101000011010011 ;
        854:  q   <=  32'b00111111000000000000000000000000 ;
        855:  q   <=  32'b00111111011100001000111110110010 ;
        856:  q   <=  32'b00111111011100001000111110110010 ;
        857:  q   <=  32'b00111111000000000000000000000000 ;
        858:  q   <=  32'b10111110001100011101000011010011 ;
        859:  q   <=  32'b10111111010001000001101101111101 ;
        860:  q   <=  32'b10111111100000000000000000000000 ;
        861:  q   <=  32'b10111111010001000001101101111101 ;
        862:  q   <=  32'b10111110001100011101000011010011 ;
        863:  q   <=  32'b00111111000000000000000000000000 ;
        864:  q   <=  32'b00111111011100001000111110110010 ;
        865:  q   <=  32'b00111111011100001000111110110010 ;
        866:  q   <=  32'b00111111000000000000000000000000 ;
        867:  q   <=  32'b10111110001100011101000011010011 ;
        868:  q   <=  32'b10111111010001000001101101111101 ;
        869:  q   <=  32'b10111111100000000000000000000000 ;
        870:  q   <=  32'b10111111010001000001101101111101 ;
        871:  q   <=  32'b10111110001100011101000011010011 ;
        872:  q   <=  32'b00111110111111111111111111111111 ;
        873:  q   <=  32'b00111111011100001000111110110010 ;
        874:  q   <=  32'b00111111011100001000111110110010 ;
        875:  q   <=  32'b00111111000000000000000000000000 ;
        876:  q   <=  32'b10111110001100011101000011010011 ;
        877:  q   <=  32'b10111111010001000001101101111101 ;
        878:  q   <=  32'b10111111100000000000000000000000 ;
        879:  q   <=  32'b10111111010001000001101101111101 ;
        880:  q   <=  32'b10111110001100011101000011010011 ;
        881:  q   <=  32'b00111110111111111111111111111111 ;
        882:  q   <=  32'b00111111011100001000111110110010 ;
        883:  q   <=  32'b00111111011011100100110110111101 ;
        884:  q   <=  32'b00111110110111100010011000000010 ;
        885:  q   <=  32'b10111110100101101110101000100110 ;
        886:  q   <=  32'b10111111010111011011001111010111 ;
        887:  q   <=  32'b10111111011110011001010011100000 ;
        888:  q   <=  32'b10111111000100000011010110111110 ;
        889:  q   <=  32'b00111110000110001001111010001001 ;
        890:  q   <=  32'b00111111010010000010011000011011 ;
        891:  q   <=  32'b00111111011111110100100010111111 ;
        892:  q   <=  32'b00111111001011100001111111001100 ;
        893:  q   <=  32'b00100101101100000111110101111101 ;
        894:  q   <=  32'b10111111001011100001111111001100 ;
        895:  q   <=  32'b10111111011111110100100010111111 ;
        896:  q   <=  32'b10111111010010000010011000011011 ;
        897:  q   <=  32'b10111110000110001001111010001001 ;
        898:  q   <=  32'b00111111000100000011010110111110 ;
        899:  q   <=  32'b00111111011110011001010011100000 ;
        900:  q   <=  32'b00111111010111011011001111010111 ;
        901:  q   <=  32'b00111110100101101110101000100110 ;
        902:  q   <=  32'b10111110110111100010011000000010 ;
        903:  q   <=  32'b10111111011011100100110110111101 ;
        904:  q   <=  32'b10111111011011100100110110111101 ;
        905:  q   <=  32'b10111110110111100010011000000010 ;
        906:  q   <=  32'b00111110100101101110101000100110 ;
        907:  q   <=  32'b00111111010111011011001111010111 ;
        908:  q   <=  32'b00111111011110011001010011100000 ;
        909:  q   <=  32'b00111111000100000011010110111110 ;
        910:  q   <=  32'b10111110000110001001111010001001 ;
        911:  q   <=  32'b10111111010010000010011000011011 ;
        912:  q   <=  32'b10111111011111110100100010111111 ;
        913:  q   <=  32'b10111111001011100001111111001100 ;
        914:  q   <=  32'b10100111010000100010111100001111 ;
        915:  q   <=  32'b00111111001011100001111111001100 ;
        916:  q   <=  32'b00111111011111110100100010111111 ;
        917:  q   <=  32'b00111111010010000010011000011011 ;
        918:  q   <=  32'b00111110000110001001111010001001 ;
        919:  q   <=  32'b10111111000100000011010110111110 ;
        920:  q   <=  32'b10111111011110011001010011100000 ;
        921:  q   <=  32'b10111111010111011011001111010111 ;
        922:  q   <=  32'b10111110100101101110101000100110 ;
        923:  q   <=  32'b00111110110111100010011000000010 ;
        924:  q   <=  32'b00111111011011100100110110111101 ;
        925:  q   <=  32'b00111111011011100100110110111101 ;
        926:  q   <=  32'b00111110110111100010011000000010 ;
        927:  q   <=  32'b10111110100101101110101000100110 ;
        928:  q   <=  32'b10111111010111011011001111010111 ;
        929:  q   <=  32'b10111111011110011001010011100000 ;
        930:  q   <=  32'b10111111000100000011010110111110 ;
        931:  q   <=  32'b00111110000110001001111010001001 ;
        932:  q   <=  32'b00111111010010000010011000011011 ;
        933:  q   <=  32'b00111111011111110100100010111111 ;
        934:  q   <=  32'b00111111001011100001111111001100 ;
        935:  q   <=  32'b10100101100011011000110010001010 ;
        936:  q   <=  32'b10111111001011100001111111001100 ;
        937:  q   <=  32'b10111111011111110100100010111111 ;
        938:  q   <=  32'b10111111010010000010011000011011 ;
        939:  q   <=  32'b10111110000110001001111010001001 ;
        940:  q   <=  32'b00111111000100000011010110111110 ;
        941:  q   <=  32'b00111111011110011001010011100000 ;
        942:  q   <=  32'b00111111010111011011001111010111 ;
        943:  q   <=  32'b00111110100101101110101000100110 ;
        944:  q   <=  32'b10111110110111100010011000000010 ;
        945:  q   <=  32'b10111111011011100100110110111101 ;
        946:  q   <=  32'b00111111011010111110010111011101 ;
        947:  q   <=  32'b00111110101110110000110111111010 ;
        948:  q   <=  32'b10111110110100101001010000111001 ;
        949:  q   <=  32'b10111111011100001000111110110010 ;
        950:  q   <=  32'b10111111011001101010010111100101 ;
        951:  q   <=  32'b10111110101000110001000010101110 ;
        952:  q   <=  32'b00111110111010011001010001110001 ;
        953:  q   <=  32'b00111111011101001010000001101011 ;
        954:  q   <=  32'b00111111011000001101001100100001 ;
        955:  q   <=  32'b00111110100010101010101110011010 ;
        956:  q   <=  32'b10111111000000000000000000000000 ;
        957:  q   <=  32'b10111111011110000001010101110010 ;
        958:  q   <=  32'b10111111010110100111000101000101 ;
        959:  q   <=  32'b10111110011000111101110010000111 ;
        960:  q   <=  32'b00111111000010101110010001001111 ;
        961:  q   <=  32'b00111111011110101110110010010101 ;
        962:  q   <=  32'b00111111010100111000010001100010 ;
        963:  q   <=  32'b00111110001100011101000011010011 ;
        964:  q   <=  32'b10111111000101010111000000111001 ;
        965:  q   <=  32'b10111111011111010010010000000100 ;
        966:  q   <=  32'b10111111010011000001000011100000 ;
        967:  q   <=  32'b10111101111111101010011111101001 ;
        968:  q   <=  32'b00111111000111111001110100000111 ;
        969:  q   <=  32'b00111111011111101011101001010110 ;
        970:  q   <=  32'b00111111010001000001101101111101 ;
        971:  q   <=  32'b00111101100110010000110000010111 ;
        972:  q   <=  32'b10111111001010010110010000111110 ;
        973:  q   <=  32'b10111111011111111010111010001000 ;
        974:  q   <=  32'b10111111001110111010100101001001 ;
        975:  q   <=  32'b10111100110011000011101101110011 ;
        976:  q   <=  32'b00111111001100101011111110100101 ;
        977:  q   <=  32'b00111111100000000000000000000000 ;
        978:  q   <=  32'b00111111001100101011111110100101 ;
        979:  q   <=  32'b10111100110011000011101101110011 ;
        980:  q   <=  32'b10111111001110111010100101001001 ;
        981:  q   <=  32'b10111111011111111010111010001000 ;
        982:  q   <=  32'b10111111001010010110010000111110 ;
        983:  q   <=  32'b00111101100110010000110000010111 ;
        984:  q   <=  32'b00111111010001000001101101111101 ;
        985:  q   <=  32'b00111111011111101011101001010110 ;
        986:  q   <=  32'b00111111000111111001110100000111 ;
        987:  q   <=  32'b10111101111111101010011111101001 ;
        988:  q   <=  32'b10111111010011000001000011100000 ;
        989:  q   <=  32'b10111111011111010010010000000100 ;
        990:  q   <=  32'b10111111000101010111000000111001 ;
        991:  q   <=  32'b00111110001100011101000011010011 ;
        992:  q   <=  32'b00111111010100111000010001100010 ;
        993:  q   <=  32'b00111111011110101110110010010101 ;
        994:  q   <=  32'b00111111000010101110010001001111 ;
        995:  q   <=  32'b10111110011000111101110010000111 ;
        996:  q   <=  32'b10111111010110100111000101000101 ;
        997:  q   <=  32'b10111111011110000001010101110010 ;
        998:  q   <=  32'b10111110111111111111111111111111 ;
        999:  q   <=  32'b00111110100010101010101110011010 ;
        1000:  q   <=  32'b00111111011000001101001100100001 ;
        1001:  q   <=  32'b00111111011101001010000001101011 ;
        1002:  q   <=  32'b00111110111010011001010001110001 ;
        1003:  q   <=  32'b10111110101000110001000010101110 ;
        1004:  q   <=  32'b10111111011001101010010111100101 ;
        1005:  q   <=  32'b10111111011100001000111110110010 ;
        1006:  q   <=  32'b10111110110100101001010000111001 ;
        1007:  q   <=  32'b00111110101110110000110111111010 ;
        1008:  q   <=  32'b00111111011010111110010111011101 ;
        1009:  q   <=  32'b00111111011010010101100001110010 ;
        1010:  q   <=  32'b00111110100101101110101000100110 ;
        1011:  q   <=  32'b10111111000001010111110011000111 ;
        1012:  q   <=  32'b10111111011111000001110001011100 ;
        1013:  q   <=  32'b10111111010010000010011000011011 ;
        1014:  q   <=  32'b10111101010011000010101100110011 ;
        1015:  q   <=  32'b00111111001101110100001100001100 ;
        1016:  q   <=  32'b00111111011111110100100010111111 ;
        1017:  q   <=  32'b00111111000110101001001011101101 ;
        1018:  q   <=  32'b10111110010010101110011011010010 ;
        1019:  q   <=  32'b10111111010111011011001111010111 ;
        1020:  q   <=  32'b10111111011100101010101101011101 ;
        1021:  q   <=  32'b10111110110001101110000011101100 ;
        1022:  q   <=  32'b00111110110111100010011000000010 ;
        1023:  q   <=  32'b00111111011101100110111010001010 ;
        1024:  q   <=  32'b00111111010101110000101111110000 ;
        1025:  q   <=  32'b00111110000110001001111010001001 ;
        1026:  q   <=  32'b10111111001001001000110110111010 ;
        1027:  q   <=  32'b10111111011111111110101110100001 ;
        1028:  q   <=  32'b10111111001011100001111111001100 ;
        1029:  q   <=  32'b00111101110010111110101000111010 ;
        1030:  q   <=  32'b00111111010011111101101100101011 ;
        1031:  q   <=  32'b00111111011110011001010011100000 ;
        1032:  q   <=  32'b00111110111101001101110110110100 ;
        1033:  q   <=  32'b10111110101011110001110101000011 ;
        1034:  q   <=  32'b10111111011011100100110110111101 ;
        1035:  q   <=  32'b10111111011000111100111010100011 ;
        1036:  q   <=  32'b10111110011111001010110111111000 ;
        1037:  q   <=  32'b00111111000100000011010110111110 ;
        1038:  q   <=  32'b00111111011111100000001101100011 ;
        1039:  q   <=  32'b00111111001111111111000110101001 ;
        1040:  q   <=  32'b10100110010100111111011101110110 ;
        1041:  q   <=  32'b10111111001111111111000110101001 ;
        1042:  q   <=  32'b10111111011111100000001101100011 ;
        1043:  q   <=  32'b10111111000100000011010110111110 ;
        1044:  q   <=  32'b00111110011111001010110111111000 ;
        1045:  q   <=  32'b00111111011000111100111010100011 ;
        1046:  q   <=  32'b00111111011011100100110110111101 ;
        1047:  q   <=  32'b00111110101011110001110101000011 ;
        1048:  q   <=  32'b10111110111101001101110110110100 ;
        1049:  q   <=  32'b10111111011110011001010011100000 ;
        1050:  q   <=  32'b10111111010011111101101100101011 ;
        1051:  q   <=  32'b10111101110010111110101000111010 ;
        1052:  q   <=  32'b00111111001011100001111111001100 ;
        1053:  q   <=  32'b00111111011111111110101110100001 ;
        1054:  q   <=  32'b00111111001001001000110110111010 ;
        1055:  q   <=  32'b10111110000110001001111010001001 ;
        1056:  q   <=  32'b10111111010101110000101111110000 ;
        1057:  q   <=  32'b10111111011101100110111010001010 ;
        1058:  q   <=  32'b10111110110111100010011000000010 ;
        1059:  q   <=  32'b00111110110001101110000011101100 ;
        1060:  q   <=  32'b00111111011100101010101101011101 ;
        1061:  q   <=  32'b00111111010111011011001111010111 ;
        1062:  q   <=  32'b00111110010010101110011011010010 ;
        1063:  q   <=  32'b10111111000110101001001011101101 ;
        1064:  q   <=  32'b10111111011111110100100010111111 ;
        1065:  q   <=  32'b10111111001101110100001100001100 ;
        1066:  q   <=  32'b00111101010011000010101100110011 ;
        1067:  q   <=  32'b00111111010010000010011000011011 ;
        1068:  q   <=  32'b00111111011111000001110001011100 ;
        1069:  q   <=  32'b00111111000001010111110011000111 ;
        1070:  q   <=  32'b10111110100101101110101000100110 ;
        1071:  q   <=  32'b10111111011010010101100001110010 ;
        1072:  q   <=  32'b00111111011001101010010111100101 ;
        1073:  q   <=  32'b00111110011000111101110010000111 ;
        1074:  q   <=  32'b10111111000111111001110100000111 ;
        1075:  q   <=  32'b10111111100000000000000000000000 ;
        1076:  q   <=  32'b10111111000111111001110100000111 ;
        1077:  q   <=  32'b00111110011000111101110010000111 ;
        1078:  q   <=  32'b00111111011001101010010111100101 ;
        1079:  q   <=  32'b00111111011001101010010111100101 ;
        1080:  q   <=  32'b00111110011000111101110010000111 ;
        1081:  q   <=  32'b10111111000111111001110100000111 ;
        1082:  q   <=  32'b10111111100000000000000000000000 ;
        1083:  q   <=  32'b10111111000111111001110100000111 ;
        1084:  q   <=  32'b00111110011000111101110010000111 ;
        1085:  q   <=  32'b00111111011001101010010111100101 ;
        1086:  q   <=  32'b00111111011001101010010111100101 ;
        1087:  q   <=  32'b00111110011000111101110010000111 ;
        1088:  q   <=  32'b10111111000111111001110100000111 ;
        1089:  q   <=  32'b10111111100000000000000000000000 ;
        1090:  q   <=  32'b10111111000111111001110100000111 ;
        1091:  q   <=  32'b00111110011000111101110010000111 ;
        1092:  q   <=  32'b00111111011001101010010111100101 ;
        1093:  q   <=  32'b00111111011001101010010111100101 ;
        1094:  q   <=  32'b00111110011000111101110010000111 ;
        1095:  q   <=  32'b10111111000111111001110100000111 ;
        1096:  q   <=  32'b10111111100000000000000000000000 ;
        1097:  q   <=  32'b10111111000111111001110100000111 ;
        1098:  q   <=  32'b00111110011000111101110010000111 ;
        1099:  q   <=  32'b00111111011001101010010111100101 ;
        1100:  q   <=  32'b00111111011001101010010111100101 ;
        1101:  q   <=  32'b00111110011000111101110010000111 ;
        1102:  q   <=  32'b10111111000111111001110100000111 ;
        1103:  q   <=  32'b10111111100000000000000000000000 ;
        1104:  q   <=  32'b10111111000111111001110100000111 ;
        1105:  q   <=  32'b00111110011000111101110010000111 ;
        1106:  q   <=  32'b00111111011001101010010111100101 ;
        1107:  q   <=  32'b00111111011001101010010111100101 ;
        1108:  q   <=  32'b00111110011000111101110010000111 ;
        1109:  q   <=  32'b10111111000111111001110100000111 ;
        1110:  q   <=  32'b10111111100000000000000000000000 ;
        1111:  q   <=  32'b10111111000111111001110100000111 ;
        1112:  q   <=  32'b00111110011000111101110010000111 ;
        1113:  q   <=  32'b00111111011001101010010111100101 ;
        1114:  q   <=  32'b00111111011001101010010111100101 ;
        1115:  q   <=  32'b00111110011000111101110010000111 ;
        1116:  q   <=  32'b10111111000111111001110100000111 ;
        1117:  q   <=  32'b10111111100000000000000000000000 ;
        1118:  q   <=  32'b10111111000111111001110100000111 ;
        1119:  q   <=  32'b00111110011000111101110010000111 ;
        1120:  q   <=  32'b00111111011001101010010111100101 ;
        1121:  q   <=  32'b00111111011001101010010111100101 ;
        1122:  q   <=  32'b00111110011000111101110010000111 ;
        1123:  q   <=  32'b10111111000111111001110100000111 ;
        1124:  q   <=  32'b10111111100000000000000000000000 ;
        1125:  q   <=  32'b10111111000111111001110100000111 ;
        1126:  q   <=  32'b00111110011000111101110010000111 ;
        1127:  q   <=  32'b00111111011001101010010111100101 ;
        1128:  q   <=  32'b00111111011001101010010111100101 ;
        1129:  q   <=  32'b00111110011000111101110010000111 ;
        1130:  q   <=  32'b10111111000111111001110100000111 ;
        1131:  q   <=  32'b10111111100000000000000000000000 ;
        1132:  q   <=  32'b10111111000111111001110100000111 ;
        1133:  q   <=  32'b00111110011000111101110010000111 ;
        1134:  q   <=  32'b00111111011001101010010111100101 ;
        1135:  q   <=  32'b00111111011000111100111010100011 ;
        1136:  q   <=  32'b00111110000110001001111010001001 ;
        1137:  q   <=  32'b10111111001101110100001100001100 ;
        1138:  q   <=  32'b10111111011111000001110001011100 ;
        1139:  q   <=  32'b10111110110111100010011000000010 ;
        1140:  q   <=  32'b00111110111101001101110110110100 ;
        1141:  q   <=  32'b00111111011111100000001101100011 ;
        1142:  q   <=  32'b00111111001011100001111111001100 ;
        1143:  q   <=  32'b10111110010010101110011011010010 ;
        1144:  q   <=  32'b10111111011010010101100001110010 ;
        1145:  q   <=  32'b10111111010111011011001111010111 ;
        1146:  q   <=  32'b10111101110010111110101000111010 ;
        1147:  q   <=  32'b00111111001111111111000110101001 ;
        1148:  q   <=  32'b00111111011110011001010011100000 ;
        1149:  q   <=  32'b00111110110001101110000011101100 ;
        1150:  q   <=  32'b10111111000001010111110011000111 ;
        1151:  q   <=  32'b10111111011111110100100010111111 ;
        1152:  q   <=  32'b10111111001001001000110110111010 ;
        1153:  q   <=  32'b00111110011111001010110111111000 ;
        1154:  q   <=  32'b00111111011011100100110110111101 ;
        1155:  q   <=  32'b00111111010101110000101111110000 ;
        1156:  q   <=  32'b00111101010011000010101100110011 ;
        1157:  q   <=  32'b10111111010010000010011000011011 ;
        1158:  q   <=  32'b10111111011101100110111010001010 ;
        1159:  q   <=  32'b10111110101011110001110101000011 ;
        1160:  q   <=  32'b00111111000100000011010110111110 ;
        1161:  q   <=  32'b00111111011111111110101110100001 ;
        1162:  q   <=  32'b00111111000110101001001011101101 ;
        1163:  q   <=  32'b10111110100101101110101000100110 ;
        1164:  q   <=  32'b10111111011100101010101101011101 ;
        1165:  q   <=  32'b10111111010011111101101100101011 ;
        1166:  q   <=  32'b10100111010100111101010100110101 ;
        1167:  q   <=  32'b00111111010011111101101100101011 ;
        1168:  q   <=  32'b00111111011100101010101101011101 ;
        1169:  q   <=  32'b00111110100101101110101000100110 ;
        1170:  q   <=  32'b10111111000110101001001011101101 ;
        1171:  q   <=  32'b10111111011111111110101110100001 ;
        1172:  q   <=  32'b10111111000100000011010110111110 ;
        1173:  q   <=  32'b00111110101011110001110101000011 ;
        1174:  q   <=  32'b00111111011101100110111010001010 ;
        1175:  q   <=  32'b00111111010010000010011000011011 ;
        1176:  q   <=  32'b10111101010011000010101100110011 ;
        1177:  q   <=  32'b10111111010101110000101111110000 ;
        1178:  q   <=  32'b10111111011011100100110110111101 ;
        1179:  q   <=  32'b10111110011111001010110111111000 ;
        1180:  q   <=  32'b00111111001001001000110110111010 ;
        1181:  q   <=  32'b00111111011111110100100010111111 ;
        1182:  q   <=  32'b00111111000001010111110011000111 ;
        1183:  q   <=  32'b10111110110001101110000011101100 ;
        1184:  q   <=  32'b10111111011110011001010011100000 ;
        1185:  q   <=  32'b10111111001111111111000110101001 ;
        1186:  q   <=  32'b00111101110010111110101000111010 ;
        1187:  q   <=  32'b00111111010111011011001111010111 ;
        1188:  q   <=  32'b00111111011010010101100001110010 ;
        1189:  q   <=  32'b00111110010010101110011011010010 ;
        1190:  q   <=  32'b10111111001011100001111111001100 ;
        1191:  q   <=  32'b10111111011111100000001101100011 ;
        1192:  q   <=  32'b10111110111101001101110110110100 ;
        1193:  q   <=  32'b00111110110111100010011000000010 ;
        1194:  q   <=  32'b00111111011111000001110001011100 ;
        1195:  q   <=  32'b00111111001101110100001100001100 ;
        1196:  q   <=  32'b10111110000110001001111010001001 ;
        1197:  q   <=  32'b10111111011000111100111010100011 ;
        1198:  q   <=  32'b00111111011000001101001100100001 ;
        1199:  q   <=  32'b00111101100110010000110000010111 ;
        1200:  q   <=  32'b10111111010011000001000011100000 ;
        1201:  q   <=  32'b10111111011100001000111110110010 ;
        1202:  q   <=  32'b10111110011000111101110010000111 ;
        1203:  q   <=  32'b00111111001100101011111110100101 ;
        1204:  q   <=  32'b00111111011110101110110010010101 ;
        1205:  q   <=  32'b00111110101110110000110111111010 ;
        1206:  q   <=  32'b10111111000101010111000000111001 ;
        1207:  q   <=  32'b10111111011111111010111010001000 ;
        1208:  q   <=  32'b10111110111111111111111111111111 ;
        1209:  q   <=  32'b00111110111010011001010001110001 ;
        1210:  q   <=  32'b00111111011111101011101001010110 ;
        1211:  q   <=  32'b00111111000111111001110100000111 ;
        1212:  q   <=  32'b10111110101000110001000010101110 ;
        1213:  q   <=  32'b10111111011110000001010101110010 ;
        1214:  q   <=  32'b10111111001110111010100101001001 ;
        1215:  q   <=  32'b00111110001100011101000011010011 ;
        1216:  q   <=  32'b00111111011010111110010111011101 ;
        1217:  q   <=  32'b00111111010100111000010001100010 ;
        1218:  q   <=  32'b10111100110011000011101101110011 ;
        1219:  q   <=  32'b10111111010110100111000101000101 ;
        1220:  q   <=  32'b10111111011001101010010111100101 ;
        1221:  q   <=  32'b10111101111111101010011111101001 ;
        1222:  q   <=  32'b00111111010001000001101101111101 ;
        1223:  q   <=  32'b00111111011101001010000001101011 ;
        1224:  q   <=  32'b00111110100010101010101110011010 ;
        1225:  q   <=  32'b10111111001010010110010000111110 ;
        1226:  q   <=  32'b10111111011111010010010000000100 ;
        1227:  q   <=  32'b10111110110100101001010000111001 ;
        1228:  q   <=  32'b00111111000010101110010001001111 ;
        1229:  q   <=  32'b00111111100000000000000000000000 ;
        1230:  q   <=  32'b00111111000010101110010001001111 ;
        1231:  q   <=  32'b10111110110100101001010000111001 ;
        1232:  q   <=  32'b10111111011111010010010000000100 ;
        1233:  q   <=  32'b10111111001010010110010000111110 ;
        1234:  q   <=  32'b00111110100010101010101110011010 ;
        1235:  q   <=  32'b00111111011101001010000001101011 ;
        1236:  q   <=  32'b00111111010001000001101101111101 ;
        1237:  q   <=  32'b10111101111111101010011111101001 ;
        1238:  q   <=  32'b10111111011001101010010111100101 ;
        1239:  q   <=  32'b10111111010110100111000101000101 ;
        1240:  q   <=  32'b10111100110011000011101101110011 ;
        1241:  q   <=  32'b00111111010100111000010001100010 ;
        1242:  q   <=  32'b00111111011010111110010111011101 ;
        1243:  q   <=  32'b00111110001100011101000011010011 ;
        1244:  q   <=  32'b10111111001110111010100101001001 ;
        1245:  q   <=  32'b10111111011110000001010101110010 ;
        1246:  q   <=  32'b10111110101000110001000010101110 ;
        1247:  q   <=  32'b00111111000111111001110100000111 ;
        1248:  q   <=  32'b00111111011111101011101001010110 ;
        1249:  q   <=  32'b00111110111010011001010001110001 ;
        1250:  q   <=  32'b10111110111111111111111111111111 ;
        1251:  q   <=  32'b10111111011111111010111010001000 ;
        1252:  q   <=  32'b10111111000101010111000000111001 ;
        1253:  q   <=  32'b00111110101110110000110111111010 ;
        1254:  q   <=  32'b00111111011110101110110010010101 ;
        1255:  q   <=  32'b00111111001100101011111110100101 ;
        1256:  q   <=  32'b10111110011000111101110010000111 ;
        1257:  q   <=  32'b10111111011100001000111110110010 ;
        1258:  q   <=  32'b10111111010011000001000011100000 ;
        1259:  q   <=  32'b00111101100110010000110000010111 ;
        1260:  q   <=  32'b00111111011000001101001100100001 ;
        1261:  q   <=  32'b00111111010111011011001111010111 ;
        1262:  q   <=  32'b00100100100011010011000100110001 ;
        1263:  q   <=  32'b10111111010111011011001111010111 ;
        1264:  q   <=  32'b10111111010111011011001111010111 ;
        1265:  q   <=  32'b10100101010100111100100111001010 ;
        1266:  q   <=  32'b00111111010111011011001111010111 ;
        1267:  q   <=  32'b00111111010111011011001111010111 ;
        1268:  q   <=  32'b00100101101100000111110101111101 ;
        1269:  q   <=  32'b10111111010111011011001111010111 ;
        1270:  q   <=  32'b10111111010111011011001111010111 ;
        1271:  q   <=  32'b10100101111101110001011000010110 ;
        1272:  q   <=  32'b00111111010111011011001111010111 ;
        1273:  q   <=  32'b00111111010111011011001111010111 ;
        1274:  q   <=  32'b00100110000111101101011101010111 ;
        1275:  q   <=  32'b10111111010111011011001111010111 ;
        1276:  q   <=  32'b10111111010111011011001111010111 ;
        1277:  q   <=  32'b10100111001100001000100011101001 ;
        1278:  q   <=  32'b00111111010111011011001111010111 ;
        1279:  q   <=  32'b00111111010111011011001111010111 ;
        1280:  q   <=  32'b10100110100011010100100000000111 ;
        1281:  q   <=  32'b10111111010111011011001111010111 ;
        1282:  q   <=  32'b10111111010111011011001111010111 ;
        1283:  q   <=  32'b10100111010000100010111100001111 ;
        1284:  q   <=  32'b00111111010111011011001111010111 ;
        1285:  q   <=  32'b00111111010111011011001111010111 ;
        1286:  q   <=  32'b10100110010100111111011101110110 ;
        1287:  q   <=  32'b10111111010111011011001111010111 ;
        1288:  q   <=  32'b10111111010111011011001111010111 ;
        1289:  q   <=  32'b10100111010100111101010100110101 ;
        1290:  q   <=  32'b00111111010111011011001111010111 ;
        1291:  q   <=  32'b00111111010111011011001111010111 ;
        1292:  q   <=  32'b00100111111011100101010000100100 ;
        1293:  q   <=  32'b10111111010111011011001111010111 ;
        1294:  q   <=  32'b10111111010111011011001111010111 ;
        1295:  q   <=  32'b00100111100011010100001001010010 ;
        1296:  q   <=  32'b00111111010111011011001111010111 ;
        1297:  q   <=  32'b00111111010111011011001111010111 ;
        1298:  q   <=  32'b10100101100011011000110010001010 ;
        1299:  q   <=  32'b10111111010111011011001111010111 ;
        1300:  q   <=  32'b10111111010111011011001111010111 ;
        1301:  q   <=  32'b10100111011101110010000110000001 ;
        1302:  q   <=  32'b00111111010111011011001111010111 ;
        1303:  q   <=  32'b00111111010111011011001111010111 ;
        1304:  q   <=  32'b00100111111111111111101001001010 ;
        1305:  q   <=  32'b10111111010111011011001111010111 ;
        1306:  q   <=  32'b10111111010111011011001111010111 ;
        1307:  q   <=  32'b00100111011101110011100001010111 ;
        1308:  q   <=  32'b00111111010111011011001111010111 ;
        1309:  q   <=  32'b00111111010111011011001111010111 ;
        1310:  q   <=  32'b00100101100011001101010111011001 ;
        1311:  q   <=  32'b10111111010111011011001111010111 ;
        1312:  q   <=  32'b10111111010111011011001111010111 ;
        1313:  q   <=  32'b10100111100011010011011011100111 ;
        1314:  q   <=  32'b00111111010111011011001111010111 ;
        1315:  q   <=  32'b00111111010111011011001111010111 ;
        1316:  q   <=  32'b00100110000011010000001110000101 ;
        1317:  q   <=  32'b10111111010111011011001111010111 ;
        1318:  q   <=  32'b10111111010111011011001111010111 ;
        1319:  q   <=  32'b10100111100101100000100111111010 ;
        1320:  q   <=  32'b00111111010111011011001111010111 ;
        1321:  q   <=  32'b00111111010111011011001111010111 ;
        1322:  q   <=  32'b10100111111001011000110001111100 ;
        1323:  q   <=  32'b10111111010111011011001111010111 ;
        1324:  q   <=  32'b00111111010110100111000101000101 ;
        1325:  q   <=  32'b10111101100110010000110000010111 ;
        1326:  q   <=  32'b10111111011010111110010111011101 ;
        1327:  q   <=  32'b10111111010001000001101101111101 ;
        1328:  q   <=  32'b00111110011000111101110010000111 ;
        1329:  q   <=  32'b00111111011110000001010101110010 ;
        1330:  q   <=  32'b00111111001010010110010000111110 ;
        1331:  q   <=  32'b10111110101110110000110111111010 ;
        1332:  q   <=  32'b10111111011111101011101001010110 ;
        1333:  q   <=  32'b10111111000010101110010001001111 ;
        1334:  q   <=  32'b00111111000000000000000000000000 ;
        1335:  q   <=  32'b00111111011111111010111010001000 ;
        1336:  q   <=  32'b00111110110100101001010000111001 ;
        1337:  q   <=  32'b10111111000111111001110100000111 ;
        1338:  q   <=  32'b10111111011110101110110010010101 ;
        1339:  q   <=  32'b10111110100010101010101110011010 ;
        1340:  q   <=  32'b00111111001110111010100101001001 ;
        1341:  q   <=  32'b00111111011100001000111110110010 ;
        1342:  q   <=  32'b00111101111111101010011111101001 ;
        1343:  q   <=  32'b10111111010100111000010001100010 ;
        1344:  q   <=  32'b10111111011000001101001100100001 ;
        1345:  q   <=  32'b00111100110011000011101101110011 ;
        1346:  q   <=  32'b00111111011001101010010111100101 ;
        1347:  q   <=  32'b00111111010011000001000011100000 ;
        1348:  q   <=  32'b10111110001100011101000011010011 ;
        1349:  q   <=  32'b10111111011101001010000001101011 ;
        1350:  q   <=  32'b10111111001100101011111110100101 ;
        1351:  q   <=  32'b00111110101000110001000010101110 ;
        1352:  q   <=  32'b00111111011111010010010000000100 ;
        1353:  q   <=  32'b00111111000101010111000000111001 ;
        1354:  q   <=  32'b10111110111010011001010001110001 ;
        1355:  q   <=  32'b10111111100000000000000000000000 ;
        1356:  q   <=  32'b10111110111010011001010001110001 ;
        1357:  q   <=  32'b00111111000101010111000000111001 ;
        1358:  q   <=  32'b00111111011111010010010000000100 ;
        1359:  q   <=  32'b00111110101000110001000010101110 ;
        1360:  q   <=  32'b10111111001100101011111110100101 ;
        1361:  q   <=  32'b10111111011101001010000001101011 ;
        1362:  q   <=  32'b10111110001100011101000011010011 ;
        1363:  q   <=  32'b00111111010011000001000011100000 ;
        1364:  q   <=  32'b00111111011001101010010111100101 ;
        1365:  q   <=  32'b00111100110011000011101101110011 ;
        1366:  q   <=  32'b10111111011000001101001100100001 ;
        1367:  q   <=  32'b10111111010100111000010001100010 ;
        1368:  q   <=  32'b00111101111111101010011111101001 ;
        1369:  q   <=  32'b00111111011100001000111110110010 ;
        1370:  q   <=  32'b00111111001110111010100101001001 ;
        1371:  q   <=  32'b10111110100010101010101110011010 ;
        1372:  q   <=  32'b10111111011110101110110010010101 ;
        1373:  q   <=  32'b10111111000111111001110100000111 ;
        1374:  q   <=  32'b00111110110100101001010000111001 ;
        1375:  q   <=  32'b00111111011111111010111010001000 ;
        1376:  q   <=  32'b00111111000000000000000000000000 ;
        1377:  q   <=  32'b10111111000010101110010001001111 ;
        1378:  q   <=  32'b10111111011111101011101001010110 ;
        1379:  q   <=  32'b10111110101110110000110111111010 ;
        1380:  q   <=  32'b00111111001010010110010000111110 ;
        1381:  q   <=  32'b00111111011110000001010101110010 ;
        1382:  q   <=  32'b00111110011000111101110010000111 ;
        1383:  q   <=  32'b10111111010001000001101101111101 ;
        1384:  q   <=  32'b10111111011010111110010111011101 ;
        1385:  q   <=  32'b10111101100110010000110000010111 ;
        1386:  q   <=  32'b00111111010110100111000101000101 ;
        1387:  q   <=  32'b00111111010101110000101111110000 ;
        1388:  q   <=  32'b10111110000110001001111010001001 ;
        1389:  q   <=  32'b10111111011101100110111010001010 ;
        1390:  q   <=  32'b10111111001001001000110110111010 ;
        1391:  q   <=  32'b00111110110111100010011000000010 ;
        1392:  q   <=  32'b00111111011111111110101110100001 ;
        1393:  q   <=  32'b00111110110001101110000011101100 ;
        1394:  q   <=  32'b10111111001011100001111111001100 ;
        1395:  q   <=  32'b10111111011100101010101101011101 ;
        1396:  q   <=  32'b10111101110010111110101000111010 ;
        1397:  q   <=  32'b00111111010111011011001111010111 ;
        1398:  q   <=  32'b00111111010011111101101100101011 ;
        1399:  q   <=  32'b10111110010010101110011011010010 ;
        1400:  q   <=  32'b10111111011110011001010011100000 ;
        1401:  q   <=  32'b10111111000110101001001011101101 ;
        1402:  q   <=  32'b00111110111101001101110110110100 ;
        1403:  q   <=  32'b00111111011111110100100010111111 ;
        1404:  q   <=  32'b00111110101011110001110101000011 ;
        1405:  q   <=  32'b10111111001101110100001100001100 ;
        1406:  q   <=  32'b10111111011011100100110110111101 ;
        1407:  q   <=  32'b10111101010011000010101100110011 ;
        1408:  q   <=  32'b00111111011000111100111010100011 ;
        1409:  q   <=  32'b00111111010010000010011000011011 ;
        1410:  q   <=  32'b10111110011111001010110111111000 ;
        1411:  q   <=  32'b10111111011111000001110001011100 ;
        1412:  q   <=  32'b10111111000100000011010110111110 ;
        1413:  q   <=  32'b00111111000001010111110011000111 ;
        1414:  q   <=  32'b00111111011111100000001101100011 ;
        1415:  q   <=  32'b00111110100101101110101000100110 ;
        1416:  q   <=  32'b10111111001111111111000110101001 ;
        1417:  q   <=  32'b10111111011010010101100001110010 ;
        1418:  q   <=  32'b00100111100011010100001001010010 ;
        1419:  q   <=  32'b00111111011010010101100001110010 ;
        1420:  q   <=  32'b00111111001111111111000110101001 ;
        1421:  q   <=  32'b10111110100101101110101000100110 ;
        1422:  q   <=  32'b10111111011111100000001101100011 ;
        1423:  q   <=  32'b10111111000001010111110011000111 ;
        1424:  q   <=  32'b00111111000100000011010110111110 ;
        1425:  q   <=  32'b00111111011111000001110001011100 ;
        1426:  q   <=  32'b00111110011111001010110111111000 ;
        1427:  q   <=  32'b10111111010010000010011000011011 ;
        1428:  q   <=  32'b10111111011000111100111010100011 ;
        1429:  q   <=  32'b00111101010011000010101100110011 ;
        1430:  q   <=  32'b00111111011011100100110110111101 ;
        1431:  q   <=  32'b00111111001101110100001100001100 ;
        1432:  q   <=  32'b10111110101011110001110101000011 ;
        1433:  q   <=  32'b10111111011111110100100010111111 ;
        1434:  q   <=  32'b10111110111101001101110110110100 ;
        1435:  q   <=  32'b00111111000110101001001011101101 ;
        1436:  q   <=  32'b00111111011110011001010011100000 ;
        1437:  q   <=  32'b00111110010010101110011011010010 ;
        1438:  q   <=  32'b10111111010011111101101100101011 ;
        1439:  q   <=  32'b10111111010111011011001111010111 ;
        1440:  q   <=  32'b00111101110010111110101000111010 ;
        1441:  q   <=  32'b00111111011100101010101101011101 ;
        1442:  q   <=  32'b00111111001011100001111111001100 ;
        1443:  q   <=  32'b10111110110001101110000011101100 ;
        1444:  q   <=  32'b10111111011111111110101110100001 ;
        1445:  q   <=  32'b10111110110111100010011000000010 ;
        1446:  q   <=  32'b00111111001001001000110110111010 ;
        1447:  q   <=  32'b00111111011101100110111010001010 ;
        1448:  q   <=  32'b00111110000110001001111010001001 ;
        1449:  q   <=  32'b10111111010101110000101111110000 ;
        1450:  q   <=  32'b00111111010100111000010001100010 ;
        1451:  q   <=  32'b10111110011000111101110010000111 ;
        1452:  q   <=  32'b10111111011111010010010000000100 ;
        1453:  q   <=  32'b10111110111111111111111111111111 ;
        1454:  q   <=  32'b00111111000111111001110100000111 ;
        1455:  q   <=  32'b00111111011101001010000001101011 ;
        1456:  q   <=  32'b00111101100110010000110000010111 ;
        1457:  q   <=  32'b10111111011001101010010111100101 ;
        1458:  q   <=  32'b10111111001110111010100101001001 ;
        1459:  q   <=  32'b00111110101110110000110111111010 ;
        1460:  q   <=  32'b00111111100000000000000000000000 ;
        1461:  q   <=  32'b00111110101110110000110111111010 ;
        1462:  q   <=  32'b10111111001110111010100101001001 ;
        1463:  q   <=  32'b10111111011001101010010111100101 ;
        1464:  q   <=  32'b00111101100110010000110000010111 ;
        1465:  q   <=  32'b00111111011101001010000001101011 ;
        1466:  q   <=  32'b00111111000111111001110100000111 ;
        1467:  q   <=  32'b10111111000000000000000000000000 ;
        1468:  q   <=  32'b10111111011111010010010000000100 ;
        1469:  q   <=  32'b10111110011000111101110010000111 ;
        1470:  q   <=  32'b00111111010100111000010001100010 ;
        1471:  q   <=  32'b00111111010100111000010001100010 ;
        1472:  q   <=  32'b10111110011000111101110010000111 ;
        1473:  q   <=  32'b10111111011111010010010000000100 ;
        1474:  q   <=  32'b10111110111111111111111111111111 ;
        1475:  q   <=  32'b00111111000111111001110100000111 ;
        1476:  q   <=  32'b00111111011101001010000001101011 ;
        1477:  q   <=  32'b00111101100110010000110000010111 ;
        1478:  q   <=  32'b10111111011001101010010111100101 ;
        1479:  q   <=  32'b10111111001110111010100101001001 ;
        1480:  q   <=  32'b00111110101110110000110111111010 ;
        1481:  q   <=  32'b00111111100000000000000000000000 ;
        1482:  q   <=  32'b00111110101110110000110111111010 ;
        1483:  q   <=  32'b10111111001110111010100101001001 ;
        1484:  q   <=  32'b10111111011001101010010111100101 ;
        1485:  q   <=  32'b00111101100110010000110000010111 ;
        1486:  q   <=  32'b00111111011101001010000001101011 ;
        1487:  q   <=  32'b00111111000111111001110100000111 ;
        1488:  q   <=  32'b10111111000000000000000000000000 ;
        1489:  q   <=  32'b10111111011111010010010000000100 ;
        1490:  q   <=  32'b10111110011000111101110010000111 ;
        1491:  q   <=  32'b00111111010100111000010001100010 ;
        1492:  q   <=  32'b00111111010100111000010001100010 ;
        1493:  q   <=  32'b10111110011000111101110010000111 ;
        1494:  q   <=  32'b10111111011111010010010000000100 ;
        1495:  q   <=  32'b10111110111111111111111111111111 ;
        1496:  q   <=  32'b00111111000111111001110100000111 ;
        1497:  q   <=  32'b00111111011101001010000001101011 ;
        1498:  q   <=  32'b00111101100110010000110000010111 ;
        1499:  q   <=  32'b10111111011001101010010111100101 ;
        1500:  q   <=  32'b10111111001110111010100101001001 ;
        1501:  q   <=  32'b00111110101110110000110111111010 ;
        1502:  q   <=  32'b00111111100000000000000000000000 ;
        1503:  q   <=  32'b00111110101110110000110111111010 ;
        1504:  q   <=  32'b10111111001110111010100101001001 ;
        1505:  q   <=  32'b10111111011001101010010111100101 ;
        1506:  q   <=  32'b00111101100110010000110000010111 ;
        1507:  q   <=  32'b00111111011101001010000001101011 ;
        1508:  q   <=  32'b00111111000111111001110100000111 ;
        1509:  q   <=  32'b10111110111111111111111111111111 ;
        1510:  q   <=  32'b10111111011111010010010000000100 ;
        1511:  q   <=  32'b10111110011000111101110010000111 ;
        1512:  q   <=  32'b00111111010100111000010001100010 ;
        1513:  q   <=  32'b00111111010011111101101100101011 ;
        1514:  q   <=  32'b10111110100101101110101000100110 ;
        1515:  q   <=  32'b10111111011111111110101110100001 ;
        1516:  q   <=  32'b10111110101011110001110101000011 ;
        1517:  q   <=  32'b00111111010010000010011000011011 ;
        1518:  q   <=  32'b00111111010101110000101111110000 ;
        1519:  q   <=  32'b10111110011111001010110111111000 ;
        1520:  q   <=  32'b10111111011111110100100010111111 ;
        1521:  q   <=  32'b10111110110001101110000011101100 ;
        1522:  q   <=  32'b00111111001111111111000110101001 ;
        1523:  q   <=  32'b00111111010111011011001111010111 ;
        1524:  q   <=  32'b10111110010010101110011011010010 ;
        1525:  q   <=  32'b10111111011111100000001101100011 ;
        1526:  q   <=  32'b10111110110111100010011000000010 ;
        1527:  q   <=  32'b00111111001101110100001100001100 ;
        1528:  q   <=  32'b00111111011000111100111010100011 ;
        1529:  q   <=  32'b10111110000110001001111010001001 ;
        1530:  q   <=  32'b10111111011111000001110001011100 ;
        1531:  q   <=  32'b10111110111101001101110110110100 ;
        1532:  q   <=  32'b00111111001011100001111111001100 ;
        1533:  q   <=  32'b00111111011010010101100001110010 ;
        1534:  q   <=  32'b10111101110010111110101000111010 ;
        1535:  q   <=  32'b10111111011110011001010011100000 ;
        1536:  q   <=  32'b10111111000001010111110011000111 ;
        1537:  q   <=  32'b00111111001001001000110110111010 ;
        1538:  q   <=  32'b00111111011011100100110110111101 ;
        1539:  q   <=  32'b10111101010011000010101100110011 ;
        1540:  q   <=  32'b10111111011101100110111010001010 ;
        1541:  q   <=  32'b10111111000100000011010110111110 ;
        1542:  q   <=  32'b00111111000110101001001011101101 ;
        1543:  q   <=  32'b00111111011100101010101101011101 ;
        1544:  q   <=  32'b10100101100011011000110010001010 ;
        1545:  q   <=  32'b10111111011100101010101101011101 ;
        1546:  q   <=  32'b10111111000110101001001011101101 ;
        1547:  q   <=  32'b00111111000100000011010110111110 ;
        1548:  q   <=  32'b00111111011101100110111010001010 ;
        1549:  q   <=  32'b00111101010011000010101100110011 ;
        1550:  q   <=  32'b10111111011011100100110110111101 ;
        1551:  q   <=  32'b10111111001001001000110110111010 ;
        1552:  q   <=  32'b00111111000001010111110011000111 ;
        1553:  q   <=  32'b00111111011110011001010011100000 ;
        1554:  q   <=  32'b00111101110010111110101000111010 ;
        1555:  q   <=  32'b10111111011010010101100001110010 ;
        1556:  q   <=  32'b10111111001011100001111111001100 ;
        1557:  q   <=  32'b00111110111101001101110110110100 ;
        1558:  q   <=  32'b00111111011111000001110001011100 ;
        1559:  q   <=  32'b00111110000110001001111010001001 ;
        1560:  q   <=  32'b10111111011000111100111010100011 ;
        1561:  q   <=  32'b10111111001101110100001100001100 ;
        1562:  q   <=  32'b00111110110111100010011000000010 ;
        1563:  q   <=  32'b00111111011111100000001101100011 ;
        1564:  q   <=  32'b00111110010010101110011011010010 ;
        1565:  q   <=  32'b10111111010111011011001111010111 ;
        1566:  q   <=  32'b10111111001111111111000110101001 ;
        1567:  q   <=  32'b00111110110001101110000011101100 ;
        1568:  q   <=  32'b00111111011111110100100010111111 ;
        1569:  q   <=  32'b00111110011111001010110111111000 ;
        1570:  q   <=  32'b10111111010101110000101111110000 ;
        1571:  q   <=  32'b10111111010010000010011000011011 ;
        1572:  q   <=  32'b00111110101011110001110101000011 ;
        1573:  q   <=  32'b00111111011111111110101110100001 ;
        1574:  q   <=  32'b00111110100101101110101000100110 ;
        1575:  q   <=  32'b10111111010011111101101100101011 ;
        1576:  q   <=  32'b00111111010011000001000011100000 ;
        1577:  q   <=  32'b10111110101110110000110111111010 ;
        1578:  q   <=  32'b10111111011111101011101001010110 ;
        1579:  q   <=  32'b10111110001100011101000011010011 ;
        1580:  q   <=  32'b00111111011001101010010111100101 ;
        1581:  q   <=  32'b00111111001010010110010000111110 ;
        1582:  q   <=  32'b10111111000010101110010001001111 ;
        1583:  q   <=  32'b10111111011101001010000001101011 ;
        1584:  q   <=  32'b00111100110011000011101101110011 ;
        1585:  q   <=  32'b00111111011110000001010101110010 ;
        1586:  q   <=  32'b00111110111111111111111111111111 ;
        1587:  q   <=  32'b10111111001100101011111110100101 ;
        1588:  q   <=  32'b10111111011000001101001100100001 ;
        1589:  q   <=  32'b00111110011000111101110010000111 ;
        1590:  q   <=  32'b00111111011111111010111010001000 ;
        1591:  q   <=  32'b00111110101000110001000010101110 ;
        1592:  q   <=  32'b10111111010100111000010001100010 ;
        1593:  q   <=  32'b10111111010001000001101101111101 ;
        1594:  q   <=  32'b00111110110100101001010000111001 ;
        1595:  q   <=  32'b00111111011111010010010000000100 ;
        1596:  q   <=  32'b00111101111111101010011111101001 ;
        1597:  q   <=  32'b10111111011010111110010111011101 ;
        1598:  q   <=  32'b10111111000111111001110100000111 ;
        1599:  q   <=  32'b00111111000101010111000000111001 ;
        1600:  q   <=  32'b00111111011100001000111110110010 ;
        1601:  q   <=  32'b10111101100110010000110000010111 ;
        1602:  q   <=  32'b10111111011110101110110010010101 ;
        1603:  q   <=  32'b10111110111010011001010001110001 ;
        1604:  q   <=  32'b00111111001110111010100101001001 ;
        1605:  q   <=  32'b00111111010110100111000101000101 ;
        1606:  q   <=  32'b10111110100010101010101110011010 ;
        1607:  q   <=  32'b10111111100000000000000000000000 ;
        1608:  q   <=  32'b10111110100010101010101110011010 ;
        1609:  q   <=  32'b00111111010110100111000101000101 ;
        1610:  q   <=  32'b00111111001110111010100101001001 ;
        1611:  q   <=  32'b10111110111010011001010001110001 ;
        1612:  q   <=  32'b10111111011110101110110010010101 ;
        1613:  q   <=  32'b10111101100110010000110000010111 ;
        1614:  q   <=  32'b00111111011100001000111110110010 ;
        1615:  q   <=  32'b00111111000101010111000000111001 ;
        1616:  q   <=  32'b10111111000111111001110100000111 ;
        1617:  q   <=  32'b10111111011010111110010111011101 ;
        1618:  q   <=  32'b00111101111111101010011111101001 ;
        1619:  q   <=  32'b00111111011111010010010000000100 ;
        1620:  q   <=  32'b00111110110100101001010000111001 ;
        1621:  q   <=  32'b10111111010001000001101101111101 ;
        1622:  q   <=  32'b10111111010100111000010001100010 ;
        1623:  q   <=  32'b00111110101000110001000010101110 ;
        1624:  q   <=  32'b00111111011111111010111010001000 ;
        1625:  q   <=  32'b00111110011000111101110010000111 ;
        1626:  q   <=  32'b10111111011000001101001100100001 ;
        1627:  q   <=  32'b10111111001100101011111110100101 ;
        1628:  q   <=  32'b00111110111111111111111111111111 ;
        1629:  q   <=  32'b00111111011110000001010101110010 ;
        1630:  q   <=  32'b00111100110011000011101101110011 ;
        1631:  q   <=  32'b10111111011101001010000001101011 ;
        1632:  q   <=  32'b10111111000010101110010001001111 ;
        1633:  q   <=  32'b00111111001010010110010000111110 ;
        1634:  q   <=  32'b00111111011001101010010111100101 ;
        1635:  q   <=  32'b10111110001100011101000011010011 ;
        1636:  q   <=  32'b10111111011111101011101001010110 ;
        1637:  q   <=  32'b10111110101110110000110111111010 ;
        1638:  q   <=  32'b00111111010011000001000011100000 ;
        1639:  q   <=  32'b00111111010010000010011000011011 ;
        1640:  q   <=  32'b10111110110111100010011000000010 ;
        1641:  q   <=  32'b10111111011110011001010011100000 ;
        1642:  q   <=  32'b10100101010100111100100111001010 ;
        1643:  q   <=  32'b00111111011110011001010011100000 ;
        1644:  q   <=  32'b00111110110111100010011000000010 ;
        1645:  q   <=  32'b10111111010010000010011000011011 ;
        1646:  q   <=  32'b10111111010010000010011000011011 ;
        1647:  q   <=  32'b00111110110111100010011000000010 ;
        1648:  q   <=  32'b00111111011110011001010011100000 ;
        1649:  q   <=  32'b00100110000111101101011101010111 ;
        1650:  q   <=  32'b10111111011110011001010011100000 ;
        1651:  q   <=  32'b10111110110111100010011000000010 ;
        1652:  q   <=  32'b00111111010010000010011000011011 ;
        1653:  q   <=  32'b00111111010010000010011000011011 ;
        1654:  q   <=  32'b10111110110111100010011000000010 ;
        1655:  q   <=  32'b10111111011110011001010011100000 ;
        1656:  q   <=  32'b10100111010000100010111100001111 ;
        1657:  q   <=  32'b00111111011110011001010011100000 ;
        1658:  q   <=  32'b00111110110111100010011000000010 ;
        1659:  q   <=  32'b10111111010010000010011000011011 ;
        1660:  q   <=  32'b10111111010010000010011000011011 ;
        1661:  q   <=  32'b00111110110111100010011000000010 ;
        1662:  q   <=  32'b00111111011110011001010011100000 ;
        1663:  q   <=  32'b00100111111011100101010000100100 ;
        1664:  q   <=  32'b10111111011110011001010011100000 ;
        1665:  q   <=  32'b10111110110111100010011000000010 ;
        1666:  q   <=  32'b00111111010010000010011000011011 ;
        1667:  q   <=  32'b00111111010010000010011000011011 ;
        1668:  q   <=  32'b10111110110111100010011000000010 ;
        1669:  q   <=  32'b10111111011110011001010011100000 ;
        1670:  q   <=  32'b10100111011101110010000110000001 ;
        1671:  q   <=  32'b00111111011110011001010011100000 ;
        1672:  q   <=  32'b00111110110111100010011000000010 ;
        1673:  q   <=  32'b10111111010010000010011000011011 ;
        1674:  q   <=  32'b10111111010010000010011000011011 ;
        1675:  q   <=  32'b00111110110111100010011000000010 ;
        1676:  q   <=  32'b00111111011110011001010011100000 ;
        1677:  q   <=  32'b00100101100011001101010111011001 ;
        1678:  q   <=  32'b10111111011110011001010011100000 ;
        1679:  q   <=  32'b10111110110111100010011000000010 ;
        1680:  q   <=  32'b00111111010010000010011000011011 ;
        1681:  q   <=  32'b00111111010010000010011000011011 ;
        1682:  q   <=  32'b10111110110111100010011000000010 ;
        1683:  q   <=  32'b10111111011110011001010011100000 ;
        1684:  q   <=  32'b10100111100101100000100111111010 ;
        1685:  q   <=  32'b00111111011110011001010011100000 ;
        1686:  q   <=  32'b00111110110111100010011000000010 ;
        1687:  q   <=  32'b10111111010010000010011000011011 ;
        1688:  q   <=  32'b10111111010010000010011000011011 ;
        1689:  q   <=  32'b00111110110111100010011000000010 ;
        1690:  q   <=  32'b00111111011110011001010011100000 ;
        1691:  q   <=  32'b00100110100011010001101001011011 ;
        1692:  q   <=  32'b10111111011110011001010011100000 ;
        1693:  q   <=  32'b10111110110111100010011000000010 ;
        1694:  q   <=  32'b00111111010010000010011000011011 ;
        1695:  q   <=  32'b00111111010010000010011000011011 ;
        1696:  q   <=  32'b10111110110111100010011000000010 ;
        1697:  q   <=  32'b10111111011110011001010011100000 ;
        1698:  q   <=  32'b10100111101100001000001100110011 ;
        1699:  q   <=  32'b00111111011110011001010011100000 ;
        1700:  q   <=  32'b00111110110111100010011000000010 ;
        1701:  q   <=  32'b10111111010010000010011000011011 ;
        1702:  q   <=  32'b00111111010001000001101101111101 ;
        1703:  q   <=  32'b10111111000000000000000000000000 ;
        1704:  q   <=  32'b10111111011100001000111110110010 ;
        1705:  q   <=  32'b00111110001100011101000011010011 ;
        1706:  q   <=  32'b00111111100000000000000000000000 ;
        1707:  q   <=  32'b00111110001100011101000011010011 ;
        1708:  q   <=  32'b10111111011100001000111110110010 ;
        1709:  q   <=  32'b10111110111111111111111111111111 ;
        1710:  q   <=  32'b00111111010001000001101101111101 ;
        1711:  q   <=  32'b00111111010001000001101101111101 ;
        1712:  q   <=  32'b10111111000000000000000000000000 ;
        1713:  q   <=  32'b10111111011100001000111110110010 ;
        1714:  q   <=  32'b00111110001100011101000011010011 ;
        1715:  q   <=  32'b00111111100000000000000000000000 ;
        1716:  q   <=  32'b00111110001100011101000011010011 ;
        1717:  q   <=  32'b10111111011100001000111110110010 ;
        1718:  q   <=  32'b10111110111111111111111111111111 ;
        1719:  q   <=  32'b00111111010001000001101101111101 ;
        1720:  q   <=  32'b00111111010001000001101101111101 ;
        1721:  q   <=  32'b10111111000000000000000000000000 ;
        1722:  q   <=  32'b10111111011100001000111110110010 ;
        1723:  q   <=  32'b00111110001100011101000011010011 ;
        1724:  q   <=  32'b00111111100000000000000000000000 ;
        1725:  q   <=  32'b00111110001100011101000011010011 ;
        1726:  q   <=  32'b10111111011100001000111110110010 ;
        1727:  q   <=  32'b10111111000000000000000000000000 ;
        1728:  q   <=  32'b00111111010001000001101101111101 ;
        1729:  q   <=  32'b00111111010001000001101101111101 ;
        1730:  q   <=  32'b10111110111111111111111111111111 ;
        1731:  q   <=  32'b10111111011100001000111110110010 ;
        1732:  q   <=  32'b00111110001100011101000011010011 ;
        1733:  q   <=  32'b00111111100000000000000000000000 ;
        1734:  q   <=  32'b00111110001100011101000011010011 ;
        1735:  q   <=  32'b10111111011100001000111110110010 ;
        1736:  q   <=  32'b10111110111111111111111111111111 ;
        1737:  q   <=  32'b00111111010001000001101101111101 ;
        1738:  q   <=  32'b00111111010001000001101101111101 ;
        1739:  q   <=  32'b10111110111111111111111111111111 ;
        1740:  q   <=  32'b10111111011100001000111110110010 ;
        1741:  q   <=  32'b00111110001100011101000011010011 ;
        1742:  q   <=  32'b00111111100000000000000000000000 ;
        1743:  q   <=  32'b00111110001100011101000011010011 ;
        1744:  q   <=  32'b10111111011100001000111110110010 ;
        1745:  q   <=  32'b10111111000000000000000000000000 ;
        1746:  q   <=  32'b00111111010001000001101101111101 ;
        1747:  q   <=  32'b00111111010001000001101101111101 ;
        1748:  q   <=  32'b10111110111111111111111111111111 ;
        1749:  q   <=  32'b10111111011100001000111110110010 ;
        1750:  q   <=  32'b00111110001100011101000011010011 ;
        1751:  q   <=  32'b00111111100000000000000000000000 ;
        1752:  q   <=  32'b00111110001100011101000011010011 ;
        1753:  q   <=  32'b10111111011100001000111110110010 ;
        1754:  q   <=  32'b10111111000000000000000000000000 ;
        1755:  q   <=  32'b00111111010001000001101101111101 ;
        1756:  q   <=  32'b00111111010001000001101101111101 ;
        1757:  q   <=  32'b10111110111111111111111111111111 ;
        1758:  q   <=  32'b10111111011100001000111110110010 ;
        1759:  q   <=  32'b00111110001100011101000011010011 ;
        1760:  q   <=  32'b00111111100000000000000000000000 ;
        1761:  q   <=  32'b00111110001100011101000011010011 ;
        1762:  q   <=  32'b10111111011100001000111110110010 ;
        1763:  q   <=  32'b10111111000000000000000000000000 ;
        1764:  q   <=  32'b00111111010001000001101101111101 ;
        1765:  q   <=  32'b00111111001111111111000110101001 ;
        1766:  q   <=  32'b10111111000100000011010110111110 ;
        1767:  q   <=  32'b10111111011000111100111010100011 ;
        1768:  q   <=  32'b00111110101011110001110101000011 ;
        1769:  q   <=  32'b00111111011110011001010011100000 ;
        1770:  q   <=  32'b10111101110010111110101000111010 ;
        1771:  q   <=  32'b10111111011111111110101110100001 ;
        1772:  q   <=  32'b10111110000110001001111010001001 ;
        1773:  q   <=  32'b00111111011101100110111010001010 ;
        1774:  q   <=  32'b00111110110001101110000011101100 ;
        1775:  q   <=  32'b10111111010111011011001111010111 ;
        1776:  q   <=  32'b10111111000110101001001011101101 ;
        1777:  q   <=  32'b00111111001101110100001100001100 ;
        1778:  q   <=  32'b00111111010010000010011000011011 ;
        1779:  q   <=  32'b10111111000001010111110011000111 ;
        1780:  q   <=  32'b10111111011010010101100001110010 ;
        1781:  q   <=  32'b00111110100101101110101000100110 ;
        1782:  q   <=  32'b00111111011111000001110001011100 ;
        1783:  q   <=  32'b10111101010011000010101100110011 ;
        1784:  q   <=  32'b10111111011111110100100010111111 ;
        1785:  q   <=  32'b10111110010010101110011011010010 ;
        1786:  q   <=  32'b00111111011100101010101101011101 ;
        1787:  q   <=  32'b00111110110111100010011000000010 ;
        1788:  q   <=  32'b10111111010101110000101111110000 ;
        1789:  q   <=  32'b10111111001001001000110110111010 ;
        1790:  q   <=  32'b00111111001011100001111111001100 ;
        1791:  q   <=  32'b00111111010011111101101100101011 ;
        1792:  q   <=  32'b10111110111101001101110110110100 ;
        1793:  q   <=  32'b10111111011011100100110110111101 ;
        1794:  q   <=  32'b00111110011111001010110111111000 ;
        1795:  q   <=  32'b00111111011111100000001101100011 ;
        1796:  q   <=  32'b00100111111111111111101001001010 ;
        1797:  q   <=  32'b10111111011111100000001101100011 ;
        1798:  q   <=  32'b10111110011111001010110111111000 ;
        1799:  q   <=  32'b00111111011011100100110110111101 ;
        1800:  q   <=  32'b00111110111101001101110110110100 ;
        1801:  q   <=  32'b10111111010011111101101100101011 ;
        1802:  q   <=  32'b10111111001011100001111111001100 ;
        1803:  q   <=  32'b00111111001001001000110110111010 ;
        1804:  q   <=  32'b00111111010101110000101111110000 ;
        1805:  q   <=  32'b10111110110111100010011000000010 ;
        1806:  q   <=  32'b10111111011100101010101101011101 ;
        1807:  q   <=  32'b00111110010010101110011011010010 ;
        1808:  q   <=  32'b00111111011111110100100010111111 ;
        1809:  q   <=  32'b00111101010011000010101100110011 ;
        1810:  q   <=  32'b10111111011111000001110001011100 ;
        1811:  q   <=  32'b10111110100101101110101000100110 ;
        1812:  q   <=  32'b00111111011010010101100001110010 ;
        1813:  q   <=  32'b00111111000001010111110011000111 ;
        1814:  q   <=  32'b10111111010010000010011000011011 ;
        1815:  q   <=  32'b10111111001101110100001100001100 ;
        1816:  q   <=  32'b00111111000110101001001011101101 ;
        1817:  q   <=  32'b00111111010111011011001111010111 ;
        1818:  q   <=  32'b10111110110001101110000011101100 ;
        1819:  q   <=  32'b10111111011101100110111010001010 ;
        1820:  q   <=  32'b00111110000110001001111010001001 ;
        1821:  q   <=  32'b00111111011111111110101110100001 ;
        1822:  q   <=  32'b00111101110010111110101000111010 ;
        1823:  q   <=  32'b10111111011110011001010011100000 ;
        1824:  q   <=  32'b10111110101011110001110101000011 ;
        1825:  q   <=  32'b00111111011000111100111010100011 ;
        1826:  q   <=  32'b00111111000100000011010110111110 ;
        1827:  q   <=  32'b10111111001111111111000110101001 ;
        1828:  q   <=  32'b00111111001110111010100101001001 ;
        1829:  q   <=  32'b10111111000111111001110100000111 ;
        1830:  q   <=  32'b10111111010100111000010001100010 ;
        1831:  q   <=  32'b00111111000000000000000000000000 ;
        1832:  q   <=  32'b00111111011001101010010111100101 ;
        1833:  q   <=  32'b10111110101110110000110111111010 ;
        1834:  q   <=  32'b10111111011101001010000001101011 ;
        1835:  q   <=  32'b00111110011000111101110010000111 ;
        1836:  q   <=  32'b00111111011111010010010000000100 ;
        1837:  q   <=  32'b10111101100110010000110000010111 ;
        1838:  q   <=  32'b10111111100000000000000000000000 ;
        1839:  q   <=  32'b10111101100110010000110000010111 ;
        1840:  q   <=  32'b00111111011111010010010000000100 ;
        1841:  q   <=  32'b00111110011000111101110010000111 ;
        1842:  q   <=  32'b10111111011101001010000001101011 ;
        1843:  q   <=  32'b10111110101110110000110111111010 ;
        1844:  q   <=  32'b00111111011001101010010111100101 ;
        1845:  q   <=  32'b00111111000000000000000000000000 ;
        1846:  q   <=  32'b10111111010100111000010001100010 ;
        1847:  q   <=  32'b10111111000111111001110100000111 ;
        1848:  q   <=  32'b00111111001110111010100101001001 ;
        1849:  q   <=  32'b00111111001110111010100101001001 ;
        1850:  q   <=  32'b10111111000111111001110100000111 ;
        1851:  q   <=  32'b10111111010100111000010001100010 ;
        1852:  q   <=  32'b00111110111111111111111111111111 ;
        1853:  q   <=  32'b00111111011001101010010111100101 ;
        1854:  q   <=  32'b10111110101110110000110111111010 ;
        1855:  q   <=  32'b10111111011101001010000001101011 ;
        1856:  q   <=  32'b00111110011000111101110010000111 ;
        1857:  q   <=  32'b00111111011111010010010000000100 ;
        1858:  q   <=  32'b10111101100110010000110000010111 ;
        1859:  q   <=  32'b10111111100000000000000000000000 ;
        1860:  q   <=  32'b10111101100110010000110000010111 ;
        1861:  q   <=  32'b00111111011111010010010000000100 ;
        1862:  q   <=  32'b00111110011000111101110010000111 ;
        1863:  q   <=  32'b10111111011101001010000001101011 ;
        1864:  q   <=  32'b10111110101110110000110111111010 ;
        1865:  q   <=  32'b00111111011001101010010111100101 ;
        1866:  q   <=  32'b00111111000000000000000000000000 ;
        1867:  q   <=  32'b10111111010100111000010001100010 ;
        1868:  q   <=  32'b10111111000111111001110100000111 ;
        1869:  q   <=  32'b00111111001110111010100101001001 ;
        1870:  q   <=  32'b00111111001110111010100101001001 ;
        1871:  q   <=  32'b10111111000111111001110100000111 ;
        1872:  q   <=  32'b10111111010100111000010001100010 ;
        1873:  q   <=  32'b00111110111111111111111111111111 ;
        1874:  q   <=  32'b00111111011001101010010111100101 ;
        1875:  q   <=  32'b10111110101110110000110111111010 ;
        1876:  q   <=  32'b10111111011101001010000001101011 ;
        1877:  q   <=  32'b00111110011000111101110010000111 ;
        1878:  q   <=  32'b00111111011111010010010000000100 ;
        1879:  q   <=  32'b10111101100110010000110000010111 ;
        1880:  q   <=  32'b10111111100000000000000000000000 ;
        1881:  q   <=  32'b10111101100110010000110000010111 ;
        1882:  q   <=  32'b00111111011111010010010000000100 ;
        1883:  q   <=  32'b00111110011000111101110010000111 ;
        1884:  q   <=  32'b10111111011101001010000001101011 ;
        1885:  q   <=  32'b10111110101110110000110111111010 ;
        1886:  q   <=  32'b00111111011001101010010111100101 ;
        1887:  q   <=  32'b00111110111111111111111111111111 ;
        1888:  q   <=  32'b10111111010100111000010001100010 ;
        1889:  q   <=  32'b10111111000111111001110100000111 ;
        1890:  q   <=  32'b00111111001110111010100101001001 ;
        1891:  q   <=  32'b00111111001101110100001100001100 ;
        1892:  q   <=  32'b10111111001011100001111111001100 ;
        1893:  q   <=  32'b10111111001111111111000110101001 ;
        1894:  q   <=  32'b00111111001001001000110110111010 ;
        1895:  q   <=  32'b00111111010010000010011000011011 ;
        1896:  q   <=  32'b10111111000110101001001011101101 ;
        1897:  q   <=  32'b10111111010011111101101100101011 ;
        1898:  q   <=  32'b00111111000100000011010110111110 ;
        1899:  q   <=  32'b00111111010101110000101111110000 ;
        1900:  q   <=  32'b10111111000001010111110011000111 ;
        1901:  q   <=  32'b10111111010111011011001111010111 ;
        1902:  q   <=  32'b00111110111101001101110110110100 ;
        1903:  q   <=  32'b00111111011000111100111010100011 ;
        1904:  q   <=  32'b10111110110111100010011000000010 ;
        1905:  q   <=  32'b10111111011010010101100001110010 ;
        1906:  q   <=  32'b00111110110001101110000011101100 ;
        1907:  q   <=  32'b00111111011011100100110110111101 ;
        1908:  q   <=  32'b10111110101011110001110101000011 ;
        1909:  q   <=  32'b10111111011100101010101101011101 ;
        1910:  q   <=  32'b00111110100101101110101000100110 ;
        1911:  q   <=  32'b00111111011101100110111010001010 ;
        1912:  q   <=  32'b10111110011111001010110111111000 ;
        1913:  q   <=  32'b10111111011110011001010011100000 ;
        1914:  q   <=  32'b00111110010010101110011011010010 ;
        1915:  q   <=  32'b00111111011111000001110001011100 ;
        1916:  q   <=  32'b10111110000110001001111010001001 ;
        1917:  q   <=  32'b10111111011111100000001101100011 ;
        1918:  q   <=  32'b00111101110010111110101000111010 ;
        1919:  q   <=  32'b00111111011111110100100010111111 ;
        1920:  q   <=  32'b10111101010011000010101100110011 ;
        1921:  q   <=  32'b10111111011111111110101110100001 ;
        1922:  q   <=  32'b00100111011101110011100001010111 ;
        1923:  q   <=  32'b00111111011111111110101110100001 ;
        1924:  q   <=  32'b00111101010011000010101100110011 ;
        1925:  q   <=  32'b10111111011111110100100010111111 ;
        1926:  q   <=  32'b10111101110010111110101000111010 ;
        1927:  q   <=  32'b00111111011111100000001101100011 ;
        1928:  q   <=  32'b00111110000110001001111010001001 ;
        1929:  q   <=  32'b10111111011111000001110001011100 ;
        1930:  q   <=  32'b10111110010010101110011011010010 ;
        1931:  q   <=  32'b00111111011110011001010011100000 ;
        1932:  q   <=  32'b00111110011111001010110111111000 ;
        1933:  q   <=  32'b10111111011101100110111010001010 ;
        1934:  q   <=  32'b10111110100101101110101000100110 ;
        1935:  q   <=  32'b00111111011100101010101101011101 ;
        1936:  q   <=  32'b00111110101011110001110101000011 ;
        1937:  q   <=  32'b10111111011011100100110110111101 ;
        1938:  q   <=  32'b10111110110001101110000011101100 ;
        1939:  q   <=  32'b00111111011010010101100001110010 ;
        1940:  q   <=  32'b00111110110111100010011000000010 ;
        1941:  q   <=  32'b10111111011000111100111010100011 ;
        1942:  q   <=  32'b10111110111101001101110110110100 ;
        1943:  q   <=  32'b00111111010111011011001111010111 ;
        1944:  q   <=  32'b00111111000001010111110011000111 ;
        1945:  q   <=  32'b10111111010101110000101111110000 ;
        1946:  q   <=  32'b10111111000100000011010110111110 ;
        1947:  q   <=  32'b00111111010011111101101100101011 ;
        1948:  q   <=  32'b00111111000110101001001011101101 ;
        1949:  q   <=  32'b10111111010010000010011000011011 ;
        1950:  q   <=  32'b10111111001001001000110110111010 ;
        1951:  q   <=  32'b00111111001111111111000110101001 ;
        1952:  q   <=  32'b00111111001011100001111111001100 ;
        1953:  q   <=  32'b10111111001101110100001100001100;
        default: q <= 0;
    endcase
end
endmodule
